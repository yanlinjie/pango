module ipsl_hmemc_ddrc_top #(
    parameter     [9:0]            TRFC_MIN                  = 10'h8c,  
    parameter     [11:0]           TREFI                     = 12'h62,  
    parameter     [5:0]            T_MRD                     = 6'h0,    
    parameter     [9:0]            T_MOD                     = 10'h0,   
    parameter                      DDR_TYPE                  = "DDR3",  
    parameter     [15:0]           MR                        = 16'h1108,
    parameter     [15:0]           EMR                       = 16'h0001,
    parameter     [15:0]           EMR2                      = 16'h0000,
    parameter     [15:0]           EMR3                      = 16'h0000,
    parameter     [6:0]            WR2PRE                    = 7'hf,
    parameter     [5:0]            T_FAW                     = 6'h10,
    parameter     [6:0]            T_RAS_MAX                 = 7'h1b,
    parameter     [5:0]            T_RAS_MIN                 = 6'hf,
    parameter     [4:0]            T_XP                      = 5'h8,
    parameter     [5:0]            RD2PRE                    = 6'h4,
    parameter     [6:0]            T_RC                      = 7'h14,
    parameter     [5:0]            WL                        = 6'h3,
    parameter     [5:0]            RL                        = 6'h5,
    parameter     [5:0]            RD2WR                     = 6'h6,
    parameter     [5:0]            WR2RD                     = 6'hd,
    parameter     [4:0]            T_RCD                     = 5'h5,
    parameter     [3:0]            T_CCD                     = 4'h4,
    parameter     [3:0]            T_RRD                     = 4'h4,
    parameter     [4:0]            T_RP                      = 5'h5,
    parameter     [3:0]            T_CKSRX                   = 4'h5,
    parameter     [3:0]            T_CKSRE                   = 4'h5,
    parameter     [5:0]            T_CKESR                   = 6'h4,
    parameter     [4:0]            T_CKE                     = 5'h3,
    parameter     [6:0]            DFI_T_RDDATA_EN           = 7'h2,
    parameter     [5:0]            DFI_TPHY_WRLAT            = 6'h2,
    parameter     [1:0]            DATA_BUS_WIDTH            = 2'b00,
    parameter                      ADDRESS_MAPPING_SEL       = 0,
    parameter                      MEM_ROW_ADDRESS           = 14,
    parameter                      MEM_COLUMN_ADDRESS        = 10,
    parameter                      MEM_BANK_ADDRESS          = 3
)(
    input                resetn,
    output               ddrc_init_done,
    input                core_clk ,
    input                ddrc_rst,
    
    input                areset_0,      
    input                aclk_0,        
                                         
    input [7:0]          awid_0,        
    input [31:0]         awaddr_0,      
    input [7:0]          awlen_0,       
    input [2:0]          awsize_0,      
    input [1:0]          awburst_0,     
    input                awlock_0,      
                                         
    input                awvalid_0,     
    output               awready_0,     
    input                awurgent_0,    
    input                awpoison_0,    
                                         
    input [127:0]        wdata_0,       
    input [15:0]         wstrb_0,       
    input                wlast_0,       
    input                wvalid_0,      
    output               wready_0,      
                                         
    output [7:0]         bid_0,         
    output [1:0]         bresp_0,       
    output               bvalid_0,      
    input                bready_0,      
                                         
    input [7:0]          arid_0,        
    input [31:0]         araddr_0,      
    input [7:0]          arlen_0,       
    input [2:0]          arsize_0,      
    input [1:0]          arburst_0,     
    input                arlock_0,      
                                         
    input                arvalid_0,     
    output               arready_0,     
    input                arpoison_0,    
                                         
    output [7:0]         rid_0,         
    output [127:0]       rdata_0,       
    output [1:0]         rresp_0,       
    output               rlast_0,       
    output               rvalid_0,      
    input                rready_0,       
    input                arurgent_0,    
    output               raq_push_0,    
    output               raq_split_0,   
    output               waq_push_0,    
    output               waq_split_0,   
                                         
    input                areset_1,      
    input                aclk_1,        
                                         
    input [7:0]          awid_1,        
    input [31:0]         awaddr_1,      
    input [7:0]          awlen_1,       
    input [2:0]          awsize_1,      
    input [1:0]          awburst_1,     
    input                awlock_1,      
                                         
    input                awvalid_1,     
    output               awready_1,     
    input                awurgent_1,    
    input                awpoison_1,    
                                         
    input [63:0]         wdata_1,       
    input [7:0]          wstrb_1,       
    input                wlast_1,       
    input                wvalid_1,      
    output               wready_1,      
                                         
    output [7:0]         bid_1,         
    output [1:0]         bresp_1,       
    output               bvalid_1,      
    input                bready_1,      
                                         
    input [7:0]          arid_1,        
    input [31:0]         araddr_1,      
    input [7:0]          arlen_1,       
    input [2:0]          arsize_1,      
    input [1:0]          arburst_1,     
    input                arlock_1,      
                                         
    input                arvalid_1,     
    output               arready_1,     
    input                arpoison_1,    
                                         
    output [7:0]         rid_1,         
    output [63:0]        rdata_1,       
    output [1:0]         rresp_1,       
    output               rlast_1,       
    output               rvalid_1,      
    input                rready_1,
                                
    input                arurgent_1,    
    output               raq_push_1,    
    output               raq_split_1,   
    output               waq_push_1,    
    output               waq_split_1,   
                                         
    input                areset_2,      
    input                aclk_2,        
                                         
    input [7:0]          awid_2,        
    input [31:0]         awaddr_2,      
    input [7:0]          awlen_2,       
    input [2:0]          awsize_2,      
    input [1:0]          awburst_2,     
    input                awlock_2,      
                                         
    input                awvalid_2,     
    output               awready_2,     
    input                awurgent_2,    
    input                awpoison_2,    
                                         
    input [63:0]         wdata_2,       
    input [7:0]          wstrb_2,       
    input                wlast_2,       
    input                wvalid_2,      
    output               wready_2,      
                                         
    output [7:0]         bid_2,         
    output [1:0]         bresp_2,       
    output               bvalid_2,      
    input                bready_2,      
                                         
    input [7:0]          arid_2,        
    input [31:0]         araddr_2,      
    input [7:0]          arlen_2,       
    input [2:0]          arsize_2,      
    input [1:0]          arburst_2,     
    input                arlock_2,      
                                         
    input                arvalid_2,     
    output               arready_2,     
    input                arpoison_2,    
                                         
    output[7:0]          rid_2,         
    output[63:0]         rdata_2,       
    output[1:0]          rresp_2,       
    output               rlast_2,       
    output               rvalid_2,      
    input                rready_2,      
                         
    input                arurgent_2,    
    output               raq_push_2,    
    output               raq_split_2,   
    output               waq_push_2,    
    output               waq_split_2,   
                                         
    input[3:0]           awqos_0,       
    input[3:0]           arqos_0,       
    input[3:0]           awqos_1,       
    input[3:0]           arqos_1,       
    input[3:0]           awqos_2,       
    input[3:0]           arqos_2,       
                                         
    input                csysreq_0,     
    output               csysack_0,     
    output               cactive_0,     
    input                csysreq_1,     
    output               csysack_1,     
    output               cactive_1,     
    input                csysreq_2,     
    output               csysack_2,     
    output               cactive_2,     
                                         
    input                csysreq_ddrc,  
    output               csysack_ddrc,  
    output               cactive_ddrc,  
    input[2:0]           pa_rmask,      
    input[2:0]           pa_wmask,
    
    input                dfi_error,            
    input[2:0]           dfi_error_info,
    input[63:0]          dfi_rddata, 
    input[3:0]           dfi_rddata_valid, 
    input                dfi_ctrlupd_ack, 
    input                dfi_phyupd_req, 
    input[1:0]           dfi_phyupd_type, 
    input                dfi_lp_ack,
    input                dfi_init_complete, 
    
    output[31:0]         dfi_address,
    output[5:0]          dfi_bank,
    output[1:0]          dfi_cas_n,
    output[1:0]          dfi_ras_n, 
    output[1:0]          dfi_we_n, 
    output[1:0]          dfi_cke,
    output[1:0]          dfi_cs,
    output[1:0]          dfi_odt,
    output[1:0]          dfi_reset_n, 
    output[63:0]         dfi_wrdata, 
    output[7:0]          dfi_wrdata_mask,
    output[3:0]          dfi_wrdata_en,
    output[3:0]          dfi_rddata_en,
    output               dfi_ctrlupd_req,
    output               dfi_dram_clk_disable, 
    output               dfi_init_start,
    output[4:0]          dfi_frequency,
    output               dfi_phyupd_ack , 
    output               dfi_lp_req,      
    output[3:0]          dfi_lp_wakeup , 

    output wire          ddrc_preset  ,
    output wire [11:0]   ddrc_paddr   ,
    output wire [31:0]   ddrc_pwdata  ,
    output wire          ddrc_pwrite  ,
    output wire          ddrc_penable ,
                    
    input                pclk,
    input                preset,
    input [11:0]         paddr,
    input [31:0]         pwdata,
    input                pwrite,
    input                penable,
    output wire          pslverr,
    input                psel,
    output wire          pready,
    output wire [31:0]   prdata 
);

  wire           ddrc_ddrc_rst    ;
  wire           ddrc_axi_reset0  ;
  wire           ddrc_axi_reset1  ;
  wire           ddrc_axi_reset2  ;
  wire           ddrc_psel    ;
  

ipsl_ddrc_reset_ctrl #(
 .TRFC_MIN            (TRFC_MIN       ),    
 .TREFI               (TREFI          ),    
 .T_MRD               (T_MRD          ),    
 .T_MOD               (T_MOD          ),    
 .DDR_TYPE            (DDR_TYPE       ),    
 .MR                  (MR             ),    
 .EMR                 (EMR            ),    
 .EMR2                (EMR2           ),    
 .EMR3                (EMR3           ),    
 .WR2PRE              (WR2PRE         ),    
 .T_FAW               (T_FAW          ),    
 .T_RAS_MAX           (T_RAS_MAX      ),    
 .T_RAS_MIN           (T_RAS_MIN      ),    
 .T_XP                (T_XP           ),    
 .RD2PRE              (RD2PRE         ),    
 .T_RC                (T_RC           ),    
 .WL                  (WL             ),    
 .RL                  (RL             ),    
 .RD2WR               (RD2WR          ),    
 .WR2RD               (WR2RD          ),    
 .T_RCD               (T_RCD          ),    
 .T_CCD               (T_CCD          ),    
 .T_RRD               (T_RRD          ),    
 .T_RP                (T_RP           ),    
 .T_CKSRX             (T_CKSRX        ),    
 .T_CKSRE             (T_CKSRE        ),    
 .T_CKESR             (T_CKESR        ),    
 .T_CKE               (T_CKE          ),    
 .DFI_T_RDDATA_EN     (DFI_T_RDDATA_EN),    
 .DFI_TPHY_WRLAT      (DFI_TPHY_WRLAT ),    
 .DATA_BUS_WIDTH      (DATA_BUS_WIDTH ),    
 .ADDRESS_MAPPING_SEL (ADDRESS_MAPPING_SEL),
 .MEM_ROW_ADDRESS     (MEM_ROW_ADDRESS    ),
 .MEM_COLUMN_ADDRESS  (MEM_COLUMN_ADDRESS ),
 .MEM_BANK_ADDRESS    (MEM_BANK_ADDRESS   ) 
)u_ipsl_ddrc_reset_ctrl (
 .pclk            (pclk           ),
 .resetn          (resetn    ),
 .user_preset     (preset    ),
 .user_pwdata     (pwdata    ),
 .user_pwrite     (pwrite    ),
 .user_penable    (penable   ),
 .user_psel       (psel      ),
 .user_paddr      (paddr     ),
 .user_ddrc_rst   (ddrc_rst  ),
 .user_axi_reset0 (areset_0),
 .user_axi_reset1 (areset_1),
 .user_axi_reset2 (areset_2),
 .ddr_init_done   (ddrc_init_done  ),
 .ddrc_rst        (ddrc_ddrc_rst    ),
 .ddrc_axi_reset0 (ddrc_axi_reset0 ),
 .ddrc_axi_reset1 (ddrc_axi_reset1 ),
 .ddrc_axi_reset2 (ddrc_axi_reset2 ),
 .ddrc_preset     (ddrc_preset     ),
 .ddrc_pwdata     (ddrc_pwdata     ),
 .ddrc_pwrite     (ddrc_pwrite     ),
 .ddrc_penable    (ddrc_penable    ),
 .ddrc_psel       (ddrc_psel       ),
 .ddrc_paddr      (ddrc_paddr      ),
 .ddrc_prdata     (prdata     ),
 .ddrc_pready     (pready     )  
);



GTP_DDRC u_ddrc(
.CORE_DDRC_CORE_CLK     (core_clk),                             
.CORE_DDRC_RST          (ddrc_ddrc_rst),                        
                        
.ARESET_0               (ddrc_axi_reset0),                   
.ACLK_0                 (aclk_0),                 
                       
.AWID_0                 (awid_0),                 
.AWADDR_0               (awaddr_0),                   
.AWLEN_0                (awlen_0),                  
.AWSIZE_0               (awsize_0),                   
.AWBURST_0              (awburst_0),                    
.AWLOCK_0               (awlock_0),                   
                        
.AWVALID_0              (awvalid_0),                    
.AWREADY_0              (awready_0),                    
.AWURGENT_0             (awurgent_0),                     
.AWPOISON_0             (awpoison_0),                     
                        
.WDATA_0                (wdata_0),                  
.WSTRB_0                (wstrb_0),                  
.WLAST_0                (wlast_0),                  
.WVALID_0               (wvalid_0),                   
.WREADY_0               (wready_0),                   
                        
.BID_0                  (bid_0),                
.BRESP_0                (bresp_0),                  
.BVALID_0               (bvalid_0),                   
.BREADY_0               (bready_0),                   
                        
.ARID_0                 (arid_0),                 
.ARADDR_0               (araddr_0),                   
.ARLEN_0                (arlen_0),                  
.ARSIZE_0               (arsize_0),                   
.ARBURST_0              (arburst_0),                    
.ARLOCK_0               (arlock_0),                   
                        
.ARVALID_0              (arvalid_0),                    
.ARREADY_0              (arready_0),                    
.ARPOISON_0             (arpoison_0),                     
                       
.RID_0                  (rid_0),                
.RDATA_0                (rdata_0),                  
.RRESP_0                (rresp_0),                  
.RLAST_0                (rlast_0),                  
.RVALID_0               (rvalid_0),                   
.RREADY_0               (rready_0),                   
.ARURGENT_0             (arurgent_0),                     
.RAQ_PUSH_0             (raq_push_0),                     
.RAQ_SPLIT_0            (raq_split_0),                                                             
.WAQ_PUSH_0             (waq_push_0),                     
.WAQ_SPLIT_0            (waq_split_0),                      
                        
.ARESET_1               (ddrc_axi_reset1),                   
.ACLK_1                 (aclk_1),                 
                       
.AWID_1                 (awid_1),                 
.AWADDR_1               (awaddr_1),                   
.AWLEN_1                (awlen_1),                  
.AWSIZE_1               (awsize_1),                   
.AWBURST_1              (awburst_1),                    
.AWLOCK_1               (awlock_1),                   
                        
.AWVALID_1              (awvalid_1),                    
.AWREADY_1              (awready_1),         
.AWURGENT_1             (awurgent_1),
.AWPOISON_1             (awpoison_1),                     
                        
.WDATA_1                (wdata_1),                  
.WSTRB_1                (wstrb_1),                  
.WLAST_1                (wlast_1),                  
.WVALID_1               (wvalid_1),                   
.WREADY_1               (wready_1),                   
                        
.BID_1                  (bid_1),                
.BRESP_1                (bresp_1),                  
.BVALID_1               (bvalid_1),                   
.BREADY_1               (bready_1),                   
                        
.ARID_1                 (arid_1),                 
.ARADDR_1               (araddr_1),                   
.ARLEN_1                (arlen_1),                  
.ARSIZE_1               (arsize_1),                   
.ARBURST_1              (arburst_1),                    
.ARLOCK_1               (arlock_1),                   
                        
.ARVALID_1              (arvalid_1),                    
.ARREADY_1              (arready_1),                    
.ARPOISON_1             (arpoison_1),                     
                       
.RID_1                  (rid_1),                
.RDATA_1                (rdata_1),                  
.RRESP_1                (rresp_1),                  
.RLAST_1                (rlast_1),                  
.RVALID_1               (rvalid_1),                   
.RREADY_1               (rready_1),                   
.ARURGENT_1             (arurgent_1),                     
.RAQ_PUSH_1             (raq_push_1),                     
.RAQ_SPLIT_1            (raq_split_1),                                                             
.WAQ_PUSH_1             (waq_push_1),                     
.WAQ_SPLIT_1            (waq_split_1),                      
                      
.ARESET_2               (ddrc_axi_reset2),                   
.ACLK_2                 (aclk_2),                 
                       
.AWID_2                 (awid_2),                 
.AWADDR_2               (awaddr_2),                   
.AWLEN_2                (awlen_2),                  
.AWSIZE_2               (awsize_2),                   
.AWBURST_2              (awburst_2),                    
.AWLOCK_2               (awlock_2),                   
                        
.AWVALID_2              (awvalid_2),                    
.AWREADY_2              (awready_2),         
.AWURGENT_2             (awurgent_2),
.AWPOISON_2             (awpoison_2),                     
                        
.WDATA_2                (wdata_2),                  
.WSTRB_2                (wstrb_2),                  
.WLAST_2                (wlast_2),                  
.WVALID_2               (wvalid_2),                   
.WREADY_2               (wready_2),                   
                        
.BID_2                  (bid_2),                
.BRESP_2                (bresp_2),                  
.BVALID_2               (bvalid_2),                   
.BREADY_2               (bready_2),                   
                        
.ARID_2                 (arid_2),                 
.ARADDR_2               (araddr_2),                   
.ARLEN_2                (arlen_2),                  
.ARSIZE_2               (arsize_2),                   
.ARBURST_2              (arburst_2),                    
.ARLOCK_2               (arlock_2),                   
                        
.ARVALID_2              (arvalid_2),                    
.ARREADY_2              (arready_2),                    
.ARPOISON_2             (arpoison_2),                     
                       
.RID_2                  (rid_2),                
.RDATA_2                (rdata_2),                  
.RRESP_2                (rresp_2),                  
.RLAST_2                (rlast_2),                  
.RVALID_2               (rvalid_2),                   
.RREADY_2               (rready_2),                   
.ARURGENT_2             (arurgent_2),                     
.RAQ_PUSH_2             (raq_push_2),                     
.RAQ_SPLIT_2            (raq_split_2),                                                             
.WAQ_PUSH_2             (waq_push_2),                     
.WAQ_SPLIT_2            (waq_split_2),     
                     
.AWQOS_0                (awqos_0),                  
.ARQOS_0                (arqos_0),                  
.AWQOS_1                (awqos_1),                  
.ARQOS_1                (arqos_1),                  
.AWQOS_2                (awqos_2),                  
.ARQOS_2                (arqos_2),                  
                       
.CSYSREQ_0              (csysreq_0),                    
.CSYSACK_0              (csysack_0),                    
.CACTIVE_0              (cactive_0),                    
.CSYSREQ_1              (csysreq_1),                    
.CSYSACK_1              (csysack_1),                    
.CACTIVE_1              (cactive_1),                    
.CSYSREQ_2              (csysreq_2),                    
.CSYSACK_2              (csysack_2),                    
.CACTIVE_2              (cactive_2),                    
                      
.CSYSREQ_DDRC           (csysreq_ddrc),                       
.CSYSACK_DDRC           (csysack_ddrc),                       
.CACTIVE_DDRC           (cactive_ddrc),                       
.PA_RMASK               (pa_rmask),                   
.PA_WMASK               (pa_wmask),                   
                    
.DFI_ADDRESS            (dfi_address),                      
.DFI_BANK               (dfi_bank),                   
.DFI_CAS_N              (dfi_cas_n),                    
.DFI_RAS_N              (dfi_ras_n),                    
.DFI_WE_N               (dfi_we_n),                   
.DFI_CKE                (dfi_cke),                  
.DFI_CS                 (dfi_cs),                 
.DFI_ODT                (dfi_odt),                  
.DFI_RESET_N            (dfi_reset_n),                      
.DFI_WRDATA             (dfi_wrdata),                     
.DFI_WRDATA_MASK        (dfi_wrdata_mask),                          
.DFI_WRDATA_EN          (dfi_wrdata_en),                        
.DFI_RDDATA             (dfi_rddata),                     
.DFI_RDDATA_EN          (dfi_rddata_en),                        
.DFI_RDDATA_VALID       (dfi_rddata_valid),                           
.DFI_CTRLUPD_ACK        (dfi_ctrlupd_ack),                                    
.DFI_CTRLUPD_REQ        (dfi_ctrlupd_req),                          
.DFI_DRAM_CLK_DISABLE   (dfi_dram_clk_disable),                                
.DFI_INIT_COMPLETE      (dfi_init_complete),                                
.DFI_INIT_START         (dfi_init_start),                         
.DFI_FREQUENCY          (dfi_frequency),                        
.DFI_PHYUPD_REQ         (dfi_phyupd_req),                            
.DFI_PHYUPD_TYPE        (dfi_phyupd_type),                            
.DFI_PHYUPD_ACK         (dfi_phyupd_ack),                            
.DFI_LP_REQ             (dfi_lp_req),                            
.DFI_LP_WAKEUP          (dfi_lp_wakeup),                            
.DFI_LP_ACK             (dfi_lp_ack),                             
.PCLK                   (pclk),               
.PRESET                 (ddrc_preset),                 
.PADDR                  (ddrc_paddr),                
.PWDATA                 (ddrc_pwdata),                 
.PWRITE                 (ddrc_pwrite),                 
.PSEL                   (ddrc_psel),               
.PENABLE                (ddrc_penable),                  
.PREADY                 (pready),                 
.PRDATA                 (prdata),                 
.PSLVERR                (pslverr)

//  .AWPOISON_INTR_2             (),
//  .ARPOISON_INTR_2             (),
//  .AWPOISON_INTR_1             (),
//  .ARPOISON_INTR_1             (),
//  .AWPOISON_INTR_0             (),
//  .ARPOISON_INTR_0             (), 
//  .RAQ_WCOUNT_0                (),
//  .RAQ_POP_0                   (),
//  .WAQ_WCOUNT_0                (),
//  .WAQ_POP_0                   (),
//  .RAQ_WCOUNT_1                (),
//  .RAQ_POP_1                   (),
//  .WAQ_WCOUNT_1                (),
//  .WAQ_POP_1                   (),
//  .RAQ_WCOUNT_2                (),
//  .RAQ_POP_2                   (),
//  .WAQ_WCOUNT_2                (),
//  .WAQ_POP_2                   (),
//  .STAT_DDRC_REG_SELFREF_TYPE (),
//  .PERF_HIF_RD_OR_WR          (),
//  .PERF_HIF_WR                (),
//  .PERF_HIF_RD                (),
//  .PERF_HIF_RMW               (),
//  .PERF_HIF_HI_PRI_RD         (),
//  .PERF_DFI_WR_DATA_CYCLES    (),
//  .PERF_DFI_RD_DATA_CYCLES    (),
//  .PERF_HPR_XACT_WHEN_CRITICAL(),
//  .PERF_LPR_XACT_WHEN_CRITICAL(),
//  .PERF_WR_XACT_WHEN_CRITICAL (),
//  .PERF_OP_IS_ACTIVATE        (),
//  .PERF_OP_IS_RD_OR_WR        (),
//  .PERF_OP_IS_RD_ACTIVATE     (),
//  .PERF_OP_IS_RD              (),
//  .PERF_OP_IS_WR              (),
//  .PERF_OP_IS_PRECHARGE       (),
//  .PERF_PRECHARGE_FOR_RDWR    (),
//  .PERF_PRECHARGE_FOR_OTHER   (),
//  .PERF_RDWR_TRANSITIONS      (),
//  .PERF_WRITE_COMBINE         (),
//  .PERF_WAR_HAZARD            (),
//  .PERF_RAW_HAZARD            (),
//  .PERF_WAW_HAZARD            (),
//  .PERF_OP_IS_ENTER_SELFREF   (),
//  .PERF_OP_IS_ENTER_POWERDOWN (),
//  .PERF_OP_IS_ENTER_DEEPPOWERDOWN (),
//  .PERF_SELFREF_MODE              (),
//  .PERF_OP_IS_REFRESH             (),
//  .PERF_OP_IS_LOAD_MODE           (),
//  .PERF_OP_IS_ZQCL                (),
//  .PERF_OP_IS_ZQCS                (),
//  .PERF_BANK                      (),
//  .PERF_HPR_REQ_WITH_NOCREDIT     (),
//  .PERF_LPR_REQ_WITH_NOCREDIT     (),
//  .LPR_CREDIT_CNT             (),
//  .HPR_CREDIT_CNT             (),
//  .WR_CREDIT_CNT              (),
//  .SCANMODE_N     (1'b1),//active low
//  .SCAN_RESET     (1'b1),
//
//  .SCAN_EN          (1'b1),
//  .RESTART_H        (),
//  .TST_DONE         (),
//  .DIAG_CLK         (1'b0),
//  .FAIL_H           (),                                           
//  .HOLD_L           (1'b0),
//  .DEBUGZ           (1'b0),
//  .DIAG_SCAN_OUT    (),
//  .TEST_H           (1'b1),
//  .BIST_CLK         (1'b0),
//  .RST_L            (1'b1)

);


endmodule