version https://git-lfs.github.com/spec/v1
oid sha256:eb9037c454c1845ac748ba8fb3505ead945658c7bf9c6ca25f0aaaafb9350555
size 915
