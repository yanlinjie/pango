version https://git-lfs.github.com/spec/v1
oid sha256:ef2f882ab93f1a255a8404dbfc9af7095a58fc86e332b927441df600caac54f1
size 1263
