version https://git-lfs.github.com/spec/v1
oid sha256:37377570718292d62f4acc3cf2e53e3a6ca4c1dd1a62bc97ea28c0ce247af27d
size 86711
