version https://git-lfs.github.com/spec/v1
oid sha256:f50a9328482e8db3d7776a5ca6db208a56c0af948dac9f08440c4c0b21861c12
size 638
