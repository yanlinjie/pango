version https://git-lfs.github.com/spec/v1
oid sha256:0a327c5a111966dc07786a16f024ca126e416bd8b042e4ef35ce8fd6396f634a
size 29868
