//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
// storage_condition module, set the storage condition, include the style: window, N-Samples
// Called by     :  debug_core
// Modification history
//
//----------------------------------------------------------------------

module ips_dbc_storage_condition_v1_3
#(
  parameter EN_WINDOWS      = 0,   //enable or disable the code simplify,0 enable;
  parameter NEW_JTAG_IF     = 1,
  parameter DATA_DEPTH = 9,            	//6~17
  parameter STOR_TYPE_CHAIN_BIT = 14,  	//{stor_type_div,stor_pos_sam}
  parameter INIT_STOR_TYPE = 0
 )
(
  input                         h_rstn ,
  input                         clk_conf ,
  input                         rst_conf ,
  input                         conf_sel ,
  input                         conf_tdi ,
  input                         shift_i ,  
  input                         clk_trig ,
  input                         rst_trig ,
  input                         trigger  ,
  input                         stor_en  ,
  output [DATA_DEPTH-1:0]       ram_wadr ,
  output                        ram_wren ,
  output                        ram_wdat0,
  output [DATA_DEPTH:0]         status,
  input                         conf_rden,
	input [4:0]                   conf_id,
	input                         conf_sel_rd,
  output                        conf_rdlast,
  output                        conf_rdata  
)/* synthesis syn_preserve = 1 */;
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity", key_keyname="SYNP15_1", key_method="rsa"
`pragma protect key_block
cvLzY2xKf6qR45ygwF2+kxmxdOElSuis1QnCGD7E9+b9o/Rggk36/stuADcEvfwAS+/26Z1lexrv
NTx+fiRVRdAxDEihrXV7oEgKoYFhneaZPM+54J5gNowv9eZrTqwbkdePBYuy24OahPOSS2Aj7yxR
kEc6vqvbTBZq7xQSuZ6ys6Rvg/R0p3Od8qmXvb9SlCmGYHuMPQ4b8lPMmyzDqKc1xoVe01gvOQ6Y
vHE1hGD4CUoVUoL5u1618YjVUAEiXxjBAcbOgkaZds9YXWdckTCuHbcdGCRsQKgXytu/4jS+xzQS
b8h6cEYtaHzld5DiPrSMehpqmDwYrg1Q1W14gg==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Pango Microsystems", key_keyname="PANGO_V1.1", key_method="rsa"
`pragma protect key_block
DMBVZabS9B+UagqUdGYfUww+Ajewx4JzLEZ+ejIugUs1fkXhuBbmFDznGMPR+Gg+jD7K7ldFFYiM
UNfd0E9UQ7wXAr8pcmP1PUkkUDz5VO5lSwFXYAMdUf92qfT1yMolAnBaMB725+1+aZC3NhmZwJgd
eXnUPscs107kATFDwkBeFamj1w5IeVqxDyJ+eJzoKI/+ig1RH4io0inhSIJCSwrg9Ub/LD4jhxmI
ha+IM/HTO4YK/DOiOhajNRLW6BYuLx+iWOz/Qvach9OP0t/EUzHtUO+sSGLZ6KM0L4STZ08FS6i3
RvmenOMQecix9D+EZ3PoFUxIAgOpBXCO63Wp5w==

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=23312)
`pragma protect data_block
l2xluHGPQyaDeHaiwZ/nCPvB1XmPLWNsHhnVORPGX+tcEmcThB/4t0uoCcMAcRnkTq2DNO/Z8wHn
G7KI48fHSUfooFE9y9gZ9IbGWyFY3XIRMbiBsmyGBzpb1qSmmH6zlt+4kYceiFdHlVQ14Em3G+JP
pGb3OdnZtS0eqHdFaSBSaQpEFrpYiNI0yovOu6144BSpz7r5VXTdh/X5DJ+88jDiLgXTuXQ8Lkbc
jurkyAmt39XfHmlRrChun+6YO61FumgpVzkLNe/BY7N6sRk6SHNXppjR1nW0V9vxEtwJ0P6I/5zu
1bt11nHZNKE3lepAsA3/F4fyKi7iJKLySIsHVvHrf2vCwweVxfxwdPYsoUtWQpYyPzXH09ieH235
JlTUyzmDG2kHLkKB6XqYzF9xRar1f1fqjBS81hOquPW4EyZjlIn7YOxACa+q6SzD1eBwNSo0wvMT
1UVmgWfMh8FOlj9PRQY6hZr/7U3zBDQkzrm00eEbOQJEtydaw19k6VGxScEhq80xiogU3DRke8Qm
jHukxVdqeDhF89pVYpuq8wNu1QFFNw4hhAyrLyp7e7O8tRqjHi/6xC52/irtpOZ0BVAGWuGSbeFz
C/5UDxzG101h2gfgNzOZn5QvLueXNxwMpqBHB4takOPelhmJB2HKw4oA6DaG2IucrW/UpTy8wzd4
gi4y2+cicsxQnXUvl/OTaWclNeLjZb23Ud/nE6djHsPJrFGJQGQ0lON3K55P3x6SG7Ppdv+acCIL
ycTftKeii/t8E8bNi8X8pJgS2jxyaOdfv3Jae/aJGjCPfshX91obmNYK2sl5kaWuLpAHyIJPBTXZ
JGRSsPOtaz9K/vJO728jWs4pSntZvVx3AjprxIVbET532wRD4rZ8rvfczWMPt3pUkwHBkeh1Xv0I
Vtg3kQT43yPrrERXlkw1RumUloZNS2i0giT/MuFnAcZ5pARiUemggY0QOxcrSw2irTNu4FyZq048
8+sh2gxBzUbpyuCpiGvA5i/SY8waxavd448RpneD09xou+9cbqtA5idIXqUc033D8VJVMtv2QaTF
oRoE/krNnokqltj3923sUlZPgE8/j93VDUELF3NTyP9hxhHZPIW5Xcl9gDbbt3AgafWutFeqe/N8
oK2qzHq14Xu539ytNadR5snC3pEyjByiPz4fB7kQnLQhArQxiy+rRzAz2VSoJgknhHVCHjGKhI5s
HDQGF50OubHqdgu9+c4I1Nv+Ic/W2+K9Hv1NBkJJ5G+G26r+Hl+L85VtBODEs1oZ3frLhAQvrl8d
8ctbDfqBfxf23yDz0kjx2c40Erc4t2RV8sLxx0yILIfmCey6AmuB85SUX7QQxqpIujL0CZ/YWQeS
KvnyfE6J3VPxfx0+IAmhWdYqkMUMbU28wpY/X9F/fvClNC1KXCW4xbN3ZFtD4KdZARVLRENd1Rx5
RwjscP01ZZsJQS0T9IbJgd+K59VW9xQxAo3wWq/FyiqrPnqH4+UVxUPPYiPVs107+rDmx1oJKSFF
qNBXKLvTJt1xC0vWIoeF+SK77xRO3GpM8sZKpLBs44sMc2p/nv+FTVwgOLo/CV3pPZtVS1Nn43dI
gqHgSl6ZaJmMTvNlIeDk3msMdfGlMYy5AxClYti4VpRqRgVv8WI981kvHweWBL7udpXfUC2Kh8wv
JzlFlf63t+8F0LgPuI0TFNF1TnHDi792JFPnLB+dtDUVRSApS7VGKvE+6iuIEYzfho+lz9wOCN4s
5eJ7V5ZXFEYcuhiNnx3mfA4YObSfYGzpoLIKTAtompE8aWS3sdzJ1/gyV9LrPMEQk3EqczTxCsHc
V03nDAv1Yiswire0vAYQ8N0CnEI/pEDaPocOnsEUZIn2vKrS40kg/PWwKuehelGLkU3mxtk55rdh
GrLbUK8Mtx2lgqc0TA6cY58g236L9PPsrrUxV4bE/cfWEG0brORzACFEctl7tZtszq5rG+pfs3Lc
kcqSrWfX7hMX+2BX5dH0AAQmpwXRPyjDZb5udu5IyjnEjKiYWuVcUXevRYwzzPN6hrRebeUGb4Pl
3aPXnKsCqZ7LxMCXLw+V4KsLQDfc45vqhTyoCL2ixFZM7wnuSFsLslWDFB/jj0DdmdcSAk7/MZ+7
sfqxaEMv+ObiJq2JhjHnHlA6FnWXJq/NMcouCf09k8Gvy2n0LPIziNCC61RY5ODMdITZBR6Cinfh
AXrXba/xqw9u65lEOeTPeFmciqNvHXH6ZLRzkgB6MZWpTJGviM6RFjAiSIuo0Fx2J2vtzb+J7l1A
R+XOKaTprsdDkPjUaXCgV7m+Po3aeL9Oyw8BdCoP1bA9tEvdxw31IKoFK1wk0kylmeZsLcQ9etLs
lor4hYQ/GYin9e4lih6ygYxvq3Ld6CIj1aMfWfFMWGOUizHe6k/7SJP6gjs3ttmdNVOS9GajoR+q
vgJt9IhBF9WY/KhLEMB5E9PdRZQbFpYUpH7Ccg0vsflqdN6ujN3IFuNcMr53XVTeWcRmmpgFsB8f
NvaCE+O7UrEyhgS/63fu4mBmrtB7j6SfAM9+1S4qef9uqQdfUJpxv3wZ82+tHXY2m16xIWFbcT1y
jXP/kIwyow8DNVXuk6axgrne7eCbT5T9E2C+Z80HoecWTq6l4/ptaMF6HhMM5QBD5leNWj/Bm65F
UzmbI+/cWuZkz6tAnDSeMxq26M5uKAiHPDjyUZQIiCX0bM6E7ng1GPUvRG/8rf07SSBei9vL7hzI
8AsAUpMp9fDukwyR9jO2yOri3DH4E0AsWEb8Kb6yseg19D54gJOELWBa+Yny9r678YYkugOp8PcJ
rP0eMOAuKRNxxgV0fJ1KeFFPnLXb3VOXVStg2DGZd2aDAqKHTMXYWTIw+RD9ma4/g6GkWKdMqxoj
dUhUdmrN1ASBZg1yiti3gOsz18GKEMRStOJvSoLYxpiq/N+OGNWgbo7EFxXLfI+LC9f1lWEOP8YM
5lw7cKwkBs/g5y+T+O8e7IABE7gC5mAMCP71nsaABKgc3tbkZkge7LkAjSwt8afi/wsjim+vZbAa
G70GwOS57ehUHf6LzeUeDiTrXs9JiibGC1LeVMPit6Tq8X5l5j2XhftwXY5KIfNlPw6Iqp6S9mIx
Q2VrdPOjdCQP/JqFRc4wiXKLy7OTJfOUh8RjNP/OcK59AtWjS0lsKE73UyTK84MxHAFAZwsZ47lg
LDhRh824hHZMX8MPAQQ2OHmiEIwyFwdNu+GtXEWQ0C/MZiPr8b1lV12Jus1LMOuetcB44vxT/fK6
Ai8tTW/AXpdoGObiVxbbFzTzUp2QeM+5TLWOqhmDa3AWgFnDcR/OEa0/HlwKwiCqSibFw0Ruzphj
lHTk72DvToqxKwYA732O4wmjUqeBqHc5sakoWEifJpn1o+hJTT4zwqoa7wUoGTqU0kCVYE7IiuYd
vE+jBpnvjPJbDNgcBm8RgkjpbwAwgJGPzlCN5y2ZA4b0dRgonqtUVJPn29hj5UO8ZXGWbyqyPvAY
nNNVPdIgant6satDYcC6jUwJFCvOaVcKwLgjVxqAgLyo/A0/64+peJ9dsOsgnj9jU41A0uwL4lGt
Dn8CyIkrcJlLQWGUtoGy8k9Ekq55uARs4jY1CfhAKdazKL4d3/TdLDCNVvwc9MzXUgpqUNTLn/Nx
z24m9Td+CAFsEzYZBUQUyYpZzuIfEVKDRRBowXzcZQPfYic9OMslTlmCskcsRoQ/5KihojO6+n22
1hy0IzqsP+KLYwOmCSORIhUFwu9UR89tWBYWWreBVgYsty+Ev7z3u2KOArMlCxxT0fiv+6xdEncq
Ilsz9QYf4nlfz3vcxc5JrW5RBGCqEwUd5HbgaiEtwxZi5PUsKbbQa6fEH0bxSHRJdg6a/Pvhft8P
8rZDTi7o0fUr5JV3WAcejo7kF6p8R3JWxgHaTAqwYJPXdzFSmFVWg6LeBndRn3HaRdqsqNmnaz+P
Im4tQjLvyPatfABgW6lO8gvQk8g/eMJTTXvmk+OakS1DKALC9iPM8vTbv6y0Ryb60nIL2h12pwhO
ARJVV2IQwLuN5RSLK0FuYozzeB4zwNCIit7eeWZiin/LdC18DTm6dgX1GukBrpNyT31khfdl4Gxz
F+JqMnTLNqIfQOZpCpX0p9j9/Y+bo15Kw4kxLC+Ov78d/vQsodEfzea9aulxR/gc+vCZn92NGq0w
YrnfjkkvucGoiqjskWBEr7T/r9xV5SjbC4XC74TvojfUyRaP33sQtXIBoIWqSllezUU/OAiTmi1K
EbeisysASZNLieIjLB6hIC9q8I+ufG0nNy1V1XExJY+oD8L2jHa8LUd/PJiT9ObCuRbrfG+UEoCO
vQP0cqVrSXDfON6pc1fSzRPyG75/raHEhIKwSohe8lalrsyIHbtoT7fxXAAkVUN6eiNJ8CaQp7jD
7BeNoXf3XkbeWPSW51O5akOopIltc+a4CNdZzgxoUfWnJhByz7DgearoqB3AC8wmw++9rWktlhK8
dhVfTb9OqIELA+FhFGnWXeRxSIwSnOYN4385zzrDG6uUor1wi6C9z0xZhQBAE5a5jOQTylNbCzU6
ohLLj29ksCsEBSbR6Rpi9WS+L2Afju2pFlMZMrPlZjGrOAL3kzfSeQgV8M7GXxsLyPJ8m8TzScpK
6GOgZHQUtuvW7UWf/jilyI2EmCYWTjNFIE8tMgZmH2bqKnd9pBqgb1c40idbr8D3GQZpNbz2qY/U
J7OYprcyCWllGo0b846ylG5duK/XuHSTLjj0MNHCdB0SckWTDIO0HJm8iVBkdLTBvbk9kAQi/xZT
vzcSADth1LnTTycO9wdI6Piqh/A78egdSJPPx0LO85iOBmt+XC5AfEoVMsm1U2251PO2qUSqH/Ei
+3Q4U25/+Yg+VHJsswu7LiGKUpnIb49xmJ8UDkGr9koBKdjPyGkUR5UJkthhp9XKzpunvUiPvkp9
j0D4k9R2w0OqGYY9PBA1OCwPghC7StJzINeyWwvZdDo82jjwcdfMrUq5/uOtLIa9OQW9PHPMIay9
nmEIxXCbOGr4d43wXIfCkfI0oZSHxaJDMLEOKv+TGlB1H+OotmG7LPvGydkuQhPRH+r8IQjH+E2k
zSpP8cpB3tV3vSZIVhkj6yRMfmAm7DIP3CZyLekTk3KKCW4pLB9fmqFvU5/SvjwPw5c63MuBq0n+
pdHrp5wsrwdxgtqcgUhj6nHjGdAJxKShS4quZihlnKrHyzmiXGba7pyJ6pNyguKj4ELlVN/Dv0Fh
Yp4Ud95sSXukapj6XsPxQNus5VC5vU5m7vw1sblSPI2wjrTfL/l0TBPLzS6WZ04ORRNd4udQUIDX
FVUyhOT7e4dbdAQC+ITRvgm1V6t+DHyJ5TTe7AizY0kTISM847SOsLK520d53oWFzw+iECh9lm30
Yktlg1GxcWNhxjRAN0OpcoqqTOg2Ds5JOUgFxJ6ptt/n2tp20gx2buqzzhrvBk2kJAdWhz+mLuVY
q9FoHfFbK9l/V22KD9CaySMZYNtGvcPmTo2Vv9Rfz7VmheDETzSuReQ2giarHubNupTJIthDXCl9
czUPzX+oCB5pi8EqivGGtHT4Amq2jyPUGDzjR/s33S/Wt3sHbTsBT/7RtQjcq0bKYHgvGsLgwNHI
cAqoRguRxVhfQ9A+ye2fgFj9OMr4+NWsBl2BrlTccP0FzIoxPUd1EYZampyePkTGKNBFoyp7lrQl
XCkyLna9/Uvi6cuuc/+EZXtYuCW7Ju9SewtvJ1iUdDBmfuZeqpo9QiZMDSyuGSTzalj8pbxV8AJ0
RtIdvhe8vbDe5Hnr1aYoOO/+uTdJR9PcxqL3HgDCIe6gmPt8vamG+cvqEAUUT69n3LCvCIJk33ZC
rZF0GZlzIuWTZV5n8qVRt0lP9rEhYPjX1PYKWU/KqDtQTf+zUjtFyQWxtQJ3nix2hQoy82GTSU/P
bC23n/ZnHKr7Tw/tzTdujl6qw7dFMusbthzWITIf+3NUFJ21tTdLEOQwPnlV83IQin6EoojFaunB
nVtmINMfM1T2v1eL4bYEp2JHrtU3E8qcEKlg9vTXaEMMugnH2KuHiLVyPCc1d9F9vMgNXCQvLM1+
asR5oOezrfZaNg9ZoTI4RnrVbR7sKsrUggf3Dibw2CsEJ63DmVfqBy5gY2lSqmmFGraEQWLqXruN
9p5YJqp6idkDr08LKUBcKnlahfFC2Gt0PodGosi25LzE92YDenf1S/XV+sd1EbrldlL0+8P6pPec
vuTj4bmPbZhakNouKyNcOis4JQi9xucO5QGDQyh+zonRIhnJO32qVw1ETz7z1uXAwzch0BE3nHmi
+ADg74pKxmWz3Jsz84xZ/PtvPt7DP3sl+1Jm/G0C94d1D/o8UX0KuamSfbw4i7G98GnGicAG/jDh
VzH198CEAybo6uqvEB8trjP1ObAr74pxFDVADDm1tNyrZp7/hZ0olMlDG9h4m2hDPF/HGuGvgdSi
eWaE4fmzCRy4aNzcPD6A/b5BG7IQscwYKF5CZR3awPml/G1OYj13B+IUBsPfZKo6ooicU2CVeUjk
G6QTGIJcJecy2HnHyo0q38RnAewRnsp8ol1CRg1pRa7msgeXNxwnaudQ8Daj+X6l4sw+DRg9UoIi
wKISanp/TcD8lqzmxfA3IVx8+dspbbmME3QMfbTIEaHpQbCuNxYZjZ47FLIwwzB+SqJkWVfbUujH
wOeMFt3BD1yKXIvoxGJUgN/mdBiYhWw5OEWB0htP5gLF3IM0M/zyap5bJ0OnDYgXyx3L9rVCsqUe
HzZIi+Oxi51n78yhgCRrhBn/3aLk+r6x86E3LaVk1UsNH3JPpZ0I3ItQ68TF9DDac0rwKBw7Qlw1
/LlK9I1Q9DJ0sdScFAFwmve3HAD1Ask1PocHGc9dhh1+MV4YyhbemxCvkBl8KPiBb8aNzakXGv5B
dfonHooPmtmag1C3jdnQSsAC5RS+CLEvWzOSGakt86Uftd41D5VgqZ0Y1FsSv7VBLitsStJfs7Pg
xsgRruJfNlILq7Rs/8KEo9OEKOCbRDyqKxm803trbP0W35TxF1xrkHSV/frZyQ87+CWCvjW1T5L9
CuBNiESFb4Gw5dkjZxQByN7lJWEQ7EXZszGZEbksdAZyq/PZ5G7ah6wlBp1ZA5IVuWolix6JtWRO
CbeRLqsmnIUdG4uSfW97Sbsjnv9SIsbrTO2p+Z9S6pjw6OO49AA1mlxH5XDjjGNOc+/4nK8krqzP
b8H1iGG0h1nL1fPZXckHNwD/ubl4a4bP+K4DBfZOwxKSgsG+DzB+vdC6tz4yN3qdUv85kOKpQo20
F4mOHZUhQRwb+u+cq7zHPFvMXSm1uVDvfI56ss9k9v4+oYKOUAtTm0AQt4hdUVB84/e9GXzmfvrn
OnuqrVMBUeyvjvyxXpV+WCDLdgw0GRs+bbcDMk20CagxIuJPap+D/hz5bCR9hjhz7vXyitdLAl2v
d0ejxBji6p8UR6/4OyvCFHLM4p3HeyacSKeNNAy7Bf+/SMhJidJbRcevDiTd53paPJbG1/IonJ14
MOKQo8UTf/xcD9emArWZ4vMtuV4hvJQzsWl74SSwbtp188BN4UtNmgvEyUJVJN07sVGVZZlSYfXC
VKlZW8kkUlkS+Gt9askwJ8KQ/6563ExfmmZJ6lHJFG2Zol3+kx0FVGX0HvkHoJK/xb9/cZzO4QJQ
UPCtd5POrjfhMlbvtA+d98UkLsr4UYI7xZNa5l4bdDJiGyQ73caLBsLuToBqFJHIQjmsuAY4ruj9
vPjZsvzcXlf4naSMhmaYFL5fKzEljo2A+OYsFu3lSDYOxyrVpKeBWz0tLZoaNWnvJJlKueQpFCnS
FTE2I2Qgo4BG/l6Hos24ximmbokWaQ7mi5DhU5Nf4XxvBkpLPW2fd0HknXmkLXoBelNE1RS87Cfe
ofRDok7pD0l0iawwuUrPzSrPqPZTHaS4dTeMDS9asw01eBlTjxPRwlkWTAM2b+T9DKZ43qq2JVS0
HBP86UO0hOBbZlgmGBKblbN5pIo5yqn9Gk+oMvMi6T1TCBmwhaxOqyMMOajUq8y8TMPw9jLmzfLf
WQzfIy03U8KWS1G7/QMnxIMdDVgQLJMrAt3LEFv9xE0TdbF+5bK/phoNleUz0niuFqtZZVp4nvnm
pTHLuJepnOMxOU10OI3VMwlRjxdavQB3S10ihRdBSeUJAFU1Ye+m/Vykr4W5YLYGQdJoj1rWmePZ
WGzp1JLhGCqqf2JRSbinYipfPrqE2GZvWkAHQUx/wNjPPxRnveTHBFhtz2dL/EB0Up1DZdENIqiX
4KMEAzchpUyZT5GQTn1WxaVngD1CRACTvK6ysIwXeGZHrQqNvSCfbzdh09LhV1P+IrzbnvKkgkX4
NVh3XNZkjcZFsGYzEH3mTsj0W5RlHmrdROiAnuDCKH9oPc7pZ/y5bDTxNrR3kKyD5FWmXbSMFkMk
0B7bVvGRkpB65ir3tZ4jZwAdek8Y4h1GcfuzqT4TbvwSguQ440ufcLLDx6yOEqNeDzknnaB7Cqst
yQozCOpWKmUwWcNu72BuRJ+EtqxIRU/caf10rLzmQOpUFIs2SR70N18XpuH2Tkzekq0CD8KfQsRf
OpbEdYbPsOUpdL4gO7wVDEZ0n2u5S0k/9b14jaY7VunKxuTFjUydFcrmHP0vaI7H0KsoFAApGDLX
PKMDvzxRbjh2ul15pJNbPJUYTigl0lPZunYQ0SnkyZV2MziNq96DyPm0f1lTvPxAY7If9Dau9DCb
i31Kf7gpsGoQIdRV8EMRR19bR518jZMIEo75I0DqBRHP7EXcb8a8EdQ40mVh7BkR7wWBv3fO5p4l
TR/KH/LPEynMM3zEdobdND+dAtyvRudda7xmMShsWhJwNmVICIZDObmxEbOaCi3H4JZp125FbkZ+
C0ffb5D/3PLEbVlX/aP7DKMkTxSfmgnbgyse0cjwNPgdLEzqoTk8duoS9BTjXKHjgA3bON76YqTe
qChVH9SFd888X1rK99e4iK3qTI0hqrd+A1Bz4/KM+57gndANIMBV8H41f4zFXfGxQ1P6qWgqpaIJ
U+VdGH196e7fk5Wza+rrrrZZi6rppZz9Lu7CtlH+7VrBY/EAfhsDDKwpBNGSHM028vWOu3Xx+F4X
yRbd+iPK/z74OkLX446JLUuQJD6jwDZaBjdJgiidFE4BGXQwb3PCjBQctL506xeYuPso/+yBeZup
T0NSUDTNXEON26/yPwwM/UYeTaDYgAr1ikxhWeQCUJu7aj+3B3M2CSM8BvOpufzGN/o504pPWqlW
WhjuOuTa0BlZ12JmDop76zNfkFtQZUi/qty2vgErjBroQAnMPWruc/2IFRgSCx06FQzgW8kVQsvg
DS06JhVVMPjFldjTN/0lLj93aoJ10Irzc/XfENYiUiQ+BrghfWO/LzgllLXiLMH9kx8HDD8219Dx
f3lrcGQYjMqxp3anVJoZH+s7b5HzaIynFElcgEhoapEJzpvuqcL6A7YVhk4EIPqkyc/F6u5fNwiy
vSYT4GvlSoLMY3liSboXLr7pobqZCxorzAXhetPrL97p8eiB28g3FeqgjAsroEwv8QlHt3awCqX5
l4DEjLiJHYDauw1ZaE93vkG5SR8E+aBD4/sA9mDdIAXuR4KltWCeAQdFSegWzR/yt/+jusqf+0gr
g/T0JZOd3l2QhC4l1Hx9QcM+1In6oi+iGerTYcLlc9ZoiPwuu/uSfrl0aWKYIe8hBLcUVyOGlEPv
dsR/5HZdtMG6kMmmjudLxYxUL31EJ3V+7No+sAaOf01x/Z+C9j9+iyPrfx2hVmzA6jZZEqs2fYgS
QOYTPL6QJdlhTu+u2dIjc28tWqdJAkpKsNh427DlrqslNwU0bYYN9+fUvn5iRU7x4/+WQfTq0LG9
cD6gm1U+dFvpT9lVjakZ6EF5ZCK/s99LATJLuid5LdXkJaz+v49DRnCE6y6QoadsbF/JFoXNbgiT
fIeKTVeVr7oOvuBwLrvGFeBL49S+2xC/5jnvRVKM7nbwabq/CnxosJDC2HhNt2DJPhN8LX3vDSff
9YKGYMcj3NkOFM7lDJGo6RpQqcLfetdtg+aVKN5zFffIlo7fi5/Bp3zoLKRDcaB5mwa8NpLBUKzM
kSnUzki5CVc8M1sb/dlNt8X35KHSDrd8FAMPrulLC+iLIK7ridUX60jHvKFdf0Sv3U9DnwZ49fJh
56DSVErCoTIS82e51onnTZ1evMPIxb8Rfv7LxIMoOJxat2iiRDkKMSYcmjzQ4BThD3hLNgJWkZVJ
vsokXzHi94AZMHPlfh1c8UnoV1fvzB++feqdShesNmYupWG4YX64QMX8EQfB5PR32M1GcC5ra2JB
IireyR1HG4vCN3ePUpDc3FSVMrlR5cjk+aJM5e3PTLWNiGuGZcZoaKZ6W1A99OJS0yKqVEq7nttp
5xmLCBJPpw8S/tpJC7MiCSgVm2u8bLMqbpFiFO1FDTit3VpgFgAxiz5JsLKN00nkkjWfCCfWiMBa
REbAVr+FEB9SOCF0Hw9BEmS9ZwImOElVzBlgtxUKjuF4bjlKc7URA84m0OEb1S5SIPwsADdeir7V
hiX5/cJ6hosHsmp7cXHXMKnAqrS4rIAvelUailUmOTslVLx7WApQlY7+XiHa8iR0aQ/epEF0vNYL
WJqU3fEGhNZc2TeGPnX/byHq7wKm+DAZoXH7gzsn9j4+4PA+vlum4hdecBnj/nrDPrJ/WU1oZYNC
7WH4pxBszspQ630WNgi/aypNmhLPlTGax3ly8BJb6NXNQSbXtsHoTVn75SuUOVyd2gq29Z+qGBq4
Km9T9wD/OD8svM50TFuR3eMxoOY2kNKe5ZyNCMAngtX4h7Uetn+EbAsWxUD612QQYWsvbIMdmP0l
kWLbC5UAxg6YxFoMcrJHRTpQDYyJ5ptyvGnKyJXaL1ZqClsAReQ0bwLuBZ01ViyytYV5rXurRgj/
1qWSwmWt9d88NA2X2MvsB6rH5v16yHl0lo6uQ20F/a+3ojQ0/9i3WWbsfVcfYm0o7tZsNCD2AqdP
KRVM4NuO3B2Z1p2NnzFtJssVy3Gr8mIrg9XwRuWp0EloXNDIBavqqeJhb/zsSfQlOo29zOSmKpNv
lgEnCpYRZl15XCr09qtMJXtD8oVNSfkJufqNLDVr7w3ZSYO+8ndkJ6d1zG7Hdk+P+8mWT5CSFnqb
KlrT84NPZHdi0+RedM2QvUU4wuuTCaIwpDCkffFDaB9paSYIb/htIfqSrxVucDeJYuveUPzNgImz
Bn8fODi67zB3sVUidwcIUD/PzYiL07Wb60wqldfL9SnkWQi2zGiueW4rtkupt8aKYAHlaJceSUoZ
ezSru8YWi8/QOyYRPrF59izFtf7gUwLI2KikALIlkWUEaF+lfnNmnhmfld5NauINnQs8/RGO1jnh
Q7WK/AVQJSCVPWaYlNjINcLPu+0QW0MLCBfwYRyd0vka/v/+BQxYQtbuY90HBV9UCbE+V1Ok+4w+
Zloolpv3If+22JWNGxgplrOL7lGMvNwR0zRfwUN960aDfz3STvVdXoA5ZUE0vNCIhokATbn3LakX
8DEIvjm+boeMAca1cEIZ8rcX2SwUwEru00qZle0q8F2+NVeyle2phhZqDYlaMSMst4R2aJzLXJsP
/hf+A++21ULZV+/OsJ1bnzEx9AIyI4gMTF+Q91zYUq6bv6wHAnFmBGJ6UF9e78r4/eHRCYYvY337
GdroZKj6Pxo4g70yTkboST0j6pBXxfRD6PODyH4RCJSIw/CFngdggxSN7sOICiNAG2v49ESbQqKf
c7QWCRTG8OXkEHnc1MAS/ZSxI/xSb/pKiMRjGiHYP6PixJXxaHsSfqV2EgmSzy7FMXL7XBEvL1Os
vmeWDBwt0f12AIvZfimoYfka3BDH/TJsddV3F86jm4gHExSoGIhUGj4jftcVZLUwaMqVvmHA+n6r
FLTYM7B1ZPBFY5aaAYSz6iXYTcvQtGzthKEh1sb9WvZ5yVfYuVRdjM8MfQJhUocdttjEILnK8Mz2
JjXdSP6+Yqz3zbXSeveOLfg6UPub+aGpLyTtJrmKCEbhuLqV4mqNRtk5BwEMrECf7w6VPgnbG/T0
TUQB6sXgeqIg9fy7PR1I4jw0VaXEeryJBE0jM3mbcJ81UrPnxRPOpihsQlBePK8i/MAP3Se0uA3c
3g8lfjNAimYhV0eGZT+N3iFVviwJ+AYcu2yyrr9zsl8tL7jV8XPnx1E6we080ldT+azdaDDFw9F4
cPaH5Wyw2RSVfXxSsaxTKBj9ytxTEPxSwoVeyq/RiTqMhgLBbNu9TV6XoXhVZFbZ2QMwGo6gHPmH
zKZ0GC8gPaERt9syhERqIiMNdxJMthpXNuCZgk/uJvMuXpBTnxDXupIS+O1Yc62dZZcrfoeLxdim
Uo5b0KxYM2+GLYsvuDfG9i9w2EaXKdzGr2tD3XjU3O5tCANpAo+JgxrDN09brUJifWDjb2Z1ufT6
wTQLUMEWBH0rRCT3fNHUL2cFnd5CxVQze9epaQbbGx1HfoekbIEL6d0bvOftPEFhmqIekDi//X2J
iRFsa5YGYJa/5F76CQGkQz264r9yhCv6fkKwbALamNrznsXHA4NgxzsEAmwo2GW5SrjtnMmFe/Gw
EiDWnxdXJ7rrxU5N6KNVumRPx4yMSE+Nw8WuczAVM+GoQF8VL2Yxt3zxy3gqOt8DFR2YujdGdono
QGNAWiwXNvmqBQICi9JxDKKRTjKsyQlNz7IYwzYtPrdnGEu2RtPbKoUpkzyM/7xCBl3EYwLtXeCS
Xgdzy3w88Ft9cfVa5Tmpz+HGRKrtSO26YjQXm5En/yMjf8J9piCYw9TPGxcajbalAQoYV3s9ftpA
GfZ0KkWWWm/ckVU9Faa+/ryFmM0YCsAEqZlOduBZADOx4SbHO63V5o99RIzr/ps/Md4fiBu4nW9/
sLftWQtMe8bKXM+E0U/pwmTjFgva1DUVe3/nzu99j/oGxPsoXmJEdwtC0+8PVdeUz6Ryb3luskmp
lLb2FkUfAy3eFtEMSPS4Z/byI5Z6HoU9pj8Xb/oC5TeHFW+nSvbee5UmTMaSjz+OubrK/ZZ4QUA3
8hzNI7PvVpL31YK6MzgchluhNfZCWDWINf6T7xAaf1ks7dy4t1/YgZeP/b48SNYbGGdINAJGKzpc
qQmTQV8MDzX9PJb9m62MLTycvzr49USS1+BkBn1AldW64BuiRE7ucQJCMeIObonpH7rqXTF6pfoU
JXWIY7FxkbTIt2HZDmnviJGpNq2HQGhvJzzGDu5iqcokA9FJZ+7eF4nr7SBXo6Q4hF4pf5Ptp9Lw
1B2jAeGh1gqVxkzpGUyfF5nl6VYMz/JvzoINSXvY6EG5bqsyrhVrs+7S+Nx4ewzSX6NQWW2wxaOL
2eGXHHaMSWIjhOn4OhCeOd1d0dsbzzuUiXANlHK4QGK9VuhlZ0w+ALCUB233AjSr3pD69mN3/XlH
85k8zdUZxG7Oi9JN1TX+ScF1I1zRO7WE3vhpcR0BWFQYthK19KIkbaSwM4bGMnJ5Q0UGPxs/UcQR
lDYkAdmoTKO3x9vQuejFY0/Eys7lTtPyiCxUr19qR7H4ryfNarZUWaXuV/TDzp6EU9lbmQEZF6YM
Gr2Yhma3TSKLoWD5kRgnLP+qPgvzahmEjet8IdYj5m2dOrx1ootkpRPOqIy9D0oHEyiNV2H2uFsb
rOQxNZBJEnN4YH2/mquGhbYyyLIeG4wbC6PVeD5a/QjHFpXod6V8Z+1bfZdCSJOyB/EvPm9CYy4/
gkWPQNrsykbrZYghAM7NAOkGoORyoIaqRMXTWKVkGGvkXRPwwoKOUpFxyZSyqS4FKB3DxjKS8LRp
XbdzIkSpkLOmLIzYMwv+4MRSkMvUdCHQ1ImPutAT2hA5TrQ1YXs+G4444SgUkuRASHbfSOGW/IiF
DfNT3S3t65axwJax6qZ4iU4r+yH1UbfF3dosyA60H1+QeZz/0CNdEVCFeAY+SSDXjjaWCIxbjJAn
ddSc14mA8wxsRZ+xHR6Ll58dsPrz5hzbNpNplZJl8mLTVc8ETMY89HnHTpmRCYBaMPsqkorffp1n
QJu8gJh3PVLYhxKTTLSLo1MDijL0zF1SWwLOuksAr+YBGBeHcXDQUAe6sl1Tih/8IQ9oVKja0XR5
OHzRBznIVe57QaFZ79f13gIZTOJouj6L34/XqDgCxnnRrxxDSpIJ7Iy3sISGtx+WBf68gArC+eFY
+0kV9vR0db0Mn1KBC1gQ/MgonELx6py2TB39mBU6g7MC0PwHQsCrvF2oRjpDhq5DNt03iLi6t68J
knEG34C+tK1SgXB7xE1dCorj3BwTUNBSBEbNlcpvspxQWWlTkFhhAzLAgpvB1Ag3QfWTyOCNxhCi
SBldGpkT0bRdTz1iv4cCeTaZ5J99jJvAdRGfPhY3RVSj0Zwmjb5mvXLAXstsYF9I7Plb0Bxl5Lm0
SPxfg5ucoTJBUeNTH+5vzAsrKa2JxwRfFzVV+VkbnMv5nAfD8JBqkEFHfmQ9frEPUTPjHrPtOCHC
5RUy2fUTx6c1wkBwX1T1HQZgDQd0D3L8hQdxQUGJlltya2ZhWXx3tXGl0DNBrdkOuYqjRXl+odI4
lM8EWwKFRYtRh+sRABoHdYXE+YKA2ag+aSCPftuJaWmAELSMBz2leCkFilJbxOb2rTpv5yjB9dWF
FOUXNH2qx6XTemWCswNKb9R24Pj2tBzn9bK5bWuYZ8qjQkwLDbw6KKC20izZxnzsE1AXfQd7+rdM
UEfU38D8ePZYVjISvUUdpgI6Lq4fCM6/SaL+1uznAhCPAT/NFpfCduMklr6LKgNQcjRBGZN0VNAa
WiiY6xBmV/D0OnV3OQ8pdIaUTwYNAc4slCeJBD6DGur9k9e6ltPhrz5V+kdSDAw/aXn11La+KuRx
t+yZYJkGKRE5mbbSPqMr7IIoI/joYdRjobKm4Qana9dIHJUEEk+QTiNnhu15iGI+7aJvAzaMRRKo
1R7nDiqXtPxoWHxYiEcLkkfeVuQBpHL0ih9WVVqmIlHsmIxXr81MWDV39xB7nTHj7QvpAtFSEUdN
3JY9cqYer9DT7C2y6TE74vK9CXdrK2IUYJ8RZD4AyI9qjeJKbbFQvtSQ3Q90+jUZbc2pAdJ5twuk
gpWVNsuPMWDc8BmVxzsT65/5Fk803OoVdMMLImb9A6D+ELe9TolREsT1GRsNvVV5hV4zrhXWHYI/
rvtMX4ieU1W3NJzERnANrdoYwLJzcmVO6WiYzx5zqZQDc38ZdmY0+zrFU36cpCIjHS2OBGAv3OeK
JtsyljwWskCAKy8TsZ8/mckY1sRGYEQ28bwBxPxgc72e+UA0eY/6Vk1OX5VfnDo/Ve28GV29nGq9
2WoMIfYzxtg8lmJ4YI+Kl5+VqSpIdbZgpTclmsvwJ5y08mJdcAAKP+yWNewrYlvhjXSXbjFt8SZs
s27LCfmdBdvfSOASMuQER5drD0nl3uEodB0zynEQpOF2kuZsBzFzakfE8w4cNLAQvljuEwiXp4/X
NYh01k0p9J1w2+DQCJlLW31ZW6E8VWhTnUu/BLvDI3q5svEjrhC/ADzg4QdyJR2bUDsZT7psAWIJ
uNv2Cio8fEGJEia5AxwAnic8fXS+g3nB/rC485SbkoL9vj1CM98cMIMYYTRZrGu9KKO8XtNVscvG
yjOJvqdr5GrIlXT46sFMEoiBBadIsWRn+LG79Y6uJ08MHQWm+cp0vqWKTNeeqSQoKWvWckpNNA37
pHJd+x7lMxhtwUEDQ89isoGWVqWjGWuenuPe0tPhqTxabYOAfLWgaq2mrpJV+dqSEuBvbZad3GQD
lE/OrrzE60r6PjBEK/buV1Vkl1J5PQE8l6fYhR2bG2Q81QR67sDC9g0hFrThcmFz7ywXfhLl0k9v
SYxta2DNFMJdhP0pha+RxQyMG81OJszJ0ZOv3lSoND2wmpoEnuoQYfwKz64p810ONZh2LVVbS1Ru
M2vMVjNp8SIOcTL1oAxSCHfkz/4fZ5aM6J2/GJi36IlnD8LoLNsgMDfH3xSIpowZhvEBJZNt3oKI
xLZKdo6FnOeCxYQTtplZa8xAMO7aDreaWXpPdgSOPnibYR1kiaSFcbbMdMvb08sTpblZ+9t1AgQw
WWGqlbrKK7D8xYJOF7V0TvAjxYeTCyrdXq7pBzSmJW3mk3cXGo4kmE5GnbjyCeoROqW2EStJjDCv
0AbIYzJPh4dGZNx9sJeDcIDqmaCfKvjC9NbN4JFmZzhnGNZyXBooFAySOdwZADyGCRcz7xoRUQ2X
m/AXjORc96iAk859hTzlRJpTF7Rti/8ygb2sxVLtFEJdRXMhvWOijDI9Qi85n8fQc/2TYeLxNmiD
y18/GmACv7d6HIt0r+oHbTJci8Fs0/kH70+SeN2tRmATdxjQlQZOtVABBrJPe3f2lDuTjTngvCtl
sLN2WiYjudapYrPemXqVA6RZLOemXrkLbIGiQUatj1ua/uLu0dXkdBKdz+Q6TbpR6ORG0pAkEN00
rs20nqwIGxQA5YVVgRLfq375vQ9dljUjJQ8DHQP9BwgLXdWLFJHOosRP8DnTJDPG646ixXL+8Rgn
hOyi88FpdAUk9ZZPKrQpnPVHvEoR5Rxy7OSe2SX9hRLtsG4xQHlqYUJbH4PGJXVySteyNH1PIMZZ
C19E+D4X1oNSEQVA5smpdKYkeNWOHnYiNMnvXJIM98ukBti+ZILM/14QwsgwLVSZoZMJU8FTJiYf
TPJ7IUI22sXnoEraKCi+jCSn7IgYQlrup6ECYXO0E6E+loRH2VW7C70K3RIRi0RgZjeGpTOTMZVt
CsR6t8z6T3f2/AE5PcjBTbzbHDfOfgidIFbQWtF28dwpA7Ym9U0DxQYkQr/7o1Zwc6RU4AdUk5eg
VDUkI/19FMCFZsuzhPx9ZqhfPgeorT27znMN/29cpLyfTbUk2b4+kn0tQweJU0J+ON5s1eWNageH
OKo7NF4I0Bco/UMX08l/XTvQs7cUelQakeJF0xUFURHb9+jNwXjL88adYTg+f9F/LWiOvvImKvKX
5XRoydM1s4Jua7QDydoj/X97NrEWJW0jM1xBNmMWl3UH6AZ0tCVZh4+65ql1wJsAmGYRXdXCmAfB
Mn7FQHsS54apIuDRBUmmuyu7KptLxCbD/+7QRWWQWWrWhhpv9rT+kTT3aCw1sDoBy2R7BhiWjBYK
yySHr2pyjzEqnMM+f5AUYuBVG5Ec0bPxwN85UNYboOPMkNwcYYrLqbs6spSuWAWKnQD1aTGderLt
o5rNZdOTAOhHqI8AdayBh8Pg1os3eeY5ZF4wiwSanNOAXYVAD+wpHm4avwsT+GX5SNaBpRmCM5oi
by2jAFHu3iybVeWAEKphnIK29eVwxp/Zh97x8YoVpqeoubyv9KY8/1s8louKBnIVBJyYwNwAg9Fz
8/MyCdl5GLWehwocW+kXE44+Lryk1k+unnu+SBLfFiUNI1W8fMRTxlhQ7rwQB2J4Wqwt0YxaPWl0
yiktWz9OM0j3WfcK50mGd13C3XufI2W+kBNcJr83AgGyIbTqBdFovd8iNDyowtP4fOiEha4SSph8
4rZvMkzgpz1+vqcXIZJZaikRLkXWRKwzaME0e+tue0yjBmtHjvhaPcULnU0tFh9uU5oONmR4h+kf
b7vYFAe6OeMunq99rQIcrhXnRlceu/Gh72H2hNlJvOaWeX4mvF849TGNnec7JG1wiFNbh8TGIqw7
/HBB9U7KHCAj/XwrJ+QhU2KHt+1Sov6sEvhsB6jr+wltjGlfy7ekVUhe8AvsctAfKG813cNm7iwE
clZ23O8LagLq96rD0EhcMzE7VX9seoIskt2MMGskweJ6LycK8DVmgzeuvSAoL5hMvJpePJ+kVEFa
jELYf2XPpBDQz8nVwBTQ4yQzgTdvY4tikU1ihRV2KWGSaCPmqIRBtGNiI/RL6sgRNAg4BbKGE82/
bm9FIUiXAjfPLHJKdd4h1okW0h+Ax4hWAQAr1PbbamLKqacSihe/lLFv0iXRpmDIpT6EK/CwAYro
uUd2X4tddEWKedZ8prp8Ox4PYrI56L/BE201rVbCLRLfHXPqc2LIIp+FmmxW1uWWgyRZqML1wzOd
fIMPEZwewLv6AE00lbB5cvADx2H6w6/hiBhIHipCfeYOCd88GFCTU8cjz1b+EDeghn8gPf/8qngF
oHUu1HyXy23sVK3wJfyHbKQMKCyDTDJF1AOSRKcMpvNwbs5IJgmyj9jtZ/1cJb1nH+T4pwm8JmLR
PMKS6oeYbWPlJZ72YegCSxoWkvCcu3TL5C3cfkrZgFjfbzDwnfi4oHMXIb5iVtontw+fdLssgqrE
hI3pXhapQCRaKc3JEvbnk6Fa8/ULuhl37jx2a88fzJPtUWjU15gKJYimSYaN8gB28t4jNMOY+Rih
WbFgToIA5kEC1ulYZHr7XpS50wS24osUxH/DwyCY9OZVFzNBQmjn6fnpPMDwxg1RWo9E1S+T4R6d
C1wsSa8euUebQAAJ/Q8PAOzK0avlJHQO3966kHP8mVkXXSswr70W13h1J5TVBk8LjScPdNC2mJQE
dhqUF+VWQEB/y3cwgCbIdsAPSvK3V/7ioMSSzHL3JVp6gPJmRlljNQKnv7ah7055jzslw+nrM67Y
Il9+PMLj6t6L7ROmtXvBTXyZYpzlHbuQ8iQOEcIaxAxTZxrF2GMhyWtfygKC83+emUIoAn2QTFil
jczmySKf6SucAqiiz2j9TK5p/U8n7PUdy/lZcUlg+rU3II9YF0Mr7K9ACn2OD1YeC2rHtKtkgelt
7QaJSNfh7VJOTCIHF8YD0Z2a5rkoMhgmWhgI/tYExvvTjaX+W+Tl4qHPLXFnC4pp3uYJqePiDBP2
O4OdcylajJ2UA2F5AS3i1d6RHxENgUhjw62Ie3Fmp/8AMT9fM3TTQAAv9KegbkupfOiXu8KlKk9Q
tQofnhmQhLE26XutcfvP/mPXTQHi8lh1OvIvSpqZmzFicuVXpqn70w4vxsUnY7CYfRONeCwKa3iF
0l6jfrHyqJhCigbRh1a3HIP1Ap+bENP/SsUMk1gN9uDXw6+1MFSFqZOhTfrxLwnjJQH01U7wOr+X
oWMLUcVtElSFiKdIrEXEZWV7Ufo8imCo+KKfwFoYCU67ieeTrfzPR/JfHQqxFZ7524Wgt11Khuw6
gfUn/3P96PqhihcwpEIY7f6qR7/6h4P+C5oAffAiDaelqVdgATiDZ+sP/wwD5yqmg3ouxHvArOQY
AblgfT6VGgnoMMn2iY9N4IcYGfgVU3pqLMlLEtsSZSK8bkenZbg48YCxq10hf6mupDL03bwnXKcX
sdzZjA9PEdXnGyqlk4nbHOJiQdiDHDRybW1q6PTyxetj23Tt58OZxoQVFidar1Hn3xKvCgk/ZUrl
/RdZfbo/vFeQ2JymB5ccIYbPj8QHM6upm6YVxaCwZRHsg8IuLwwTc7luiXRCoDGlDXFKp1JJOcpU
arAX2N1Kxb0p+EXzdMXyBc6xAFmDh5AJOSeKqONrDEAUrXBkmQ/V3Sp6d7KaHMqAGnsHbufkiUj5
SVV/x4HxEnZZsXhohISvYu2EhviVH0GQ69HyJhB5a7P4KV+izFkw5TGViKm5QQfsQ1tmcQ6iAbqZ
YEKIMZ4dLrtfyAW+u/7tO9PwKoViIkPUtzGgEk56+9UhfHa7zmIJ/hDaZW/9QeAzEgbu5TMnOuUC
EwxYZKJF63CkFnwAhXLW4+tQmK+DjtVMNS+yBThLAD0N8NyZR5OELZodtTz2HjRxksKp+30dfqW4
9shBd/uG1CA+/oVG1YuNyJVEdxyyvxl28Z2vQHir/QDs7VrGSyl7IzaulHiQU5djF+z3RgMsj5Dp
IHJtYIZxmNeu/IEXTQUvQN5JrVKLouw7sgu+FXofPvvIdSrP/JgHDA0IigoRzE+uSl30WyIdtWv4
dLUlK8wza5AtaSq1BKVbQ12N1EOvUiHhIhRkEZhg1RnATSY1oUHpRExoqjUWinzwnYh6bRaF5Uz1
IqDkO4tIMa9/l69TzRJ/nr+NF+02+ihTWlx2UDoBdo10L+Y2hyy+MZhdy1DbifyEUr+lEhwpzF5h
b7MpsjAFtDcLfBJsEp8Y3IkgnLINVd9E9Qm01WRmspkqugiHCHe5wb8wgcI4QXz6+HrUXDxpcCOe
hUEUcF78qhmLLj7tl6+NCO6+aptunkACNCf5aV2yJG9IqFTtr9bHQyp4eGKGhR4k446uOzNz2pav
AqpMjPysxYomh355qrOcE9sOUKrfsY8doPHFrU5lmxt+PfZypJCKeUDa0nEMA04szUuM1Uc48njc
X+rxjBYhtI1b/G9aVYqZQD5CJQpsW1YS9T5QFI9VzSalU0geHfRrTMshZsHU37+CpJgu+1rcyIux
5l5BS2rkcaHk+Cu8zp9m4KgZruredc/JUi4+N+YDeaClyefrEXB1D7tLxVICz6B3eXs3H2QA3hX7
ErVwRYnGh6XmDEpA/AdDZT8lve0WMu3FlrwZnX/SVE91PWGVfaWgezk+H/epyL6s4qn4glhMxSDN
2stJW2K4btd2DoBl7FDXIfbpd/wyRSKoCTWku0XvXZK9kO24u4rx5swWSr59erxXC71G5VM9xdC8
QhFZtYJHFDY1O0PEe8GAulvuXBT3DfTngyv53yei2Hp9ROfbWbJ07m6SuzY1Cggx8pQa9t+PtiAL
/bo5ECeU7jXqcxy+GoQ1w5AM1Wne7acojNl2OKIxXQ9m/e4h/V7deNgn53z7ekBFTR7du0LBatSq
7j7/RBn5E2s/kjUDPvWYvrvQEpZI2x5+mGdpaQS7QjNjtFBdWAV1m+urBU5RaRa7qFDp39qhtKLG
URCZItpap4CGNy/zsy4OI2z1+u7C17Ym1fmhtUv4AUtDMqeobTQsOhDXbr/yyC/kOvCGbqF/bHX/
ctGQW08Vf9Ab7DDLS0Eh/+CvXv7rGuFgE+mtwEpE9rLYaMrongOvzjq19S61kWSPUb8lAptHBQzO
9u+UmnpcsxxymRDNu/aMhAcHGWNaslZoZGzOJrO9smD4a1v1l3N1mV3tCAqg1l6A0fMn9aUUjZvp
6yFjsHDz/ZzK8JwdfcLGuTU/xuv49Oui7540JRDIFT1bOsO3DwLyvUgE4OpY60SyI+nPK1C/CTtH
s2eWQu3iIo2V105EkuDI6rhKtSpSn6H+0I0oD+aHzU7L+woLuMHTqpx/nn+PWqtPHWBCuIXPk/MS
tb6w900sM7PFU0+qZINmM/ZfBBcjAvxBz11XBHMGk06/sPdrNOM5Dp3x32TR+iGHjvhdgyXa7RSF
G93dtN9wUHiknBOdvs4uaYhPKRQdXg3OyAZI2OeqrFBc/4MR4UD9JPOJV1+yN3NfrRf7lSWla1lz
5y2e1Izd19p/4N5WtXk7ijgQC0ZWTPVeEaW6wRlUN/GFwuSsLwCWARODhPaUNR6oQ4pw6BwpSytt
Bo2PfXwhPCSScZA6Nu++pAATB/AqOGUZmqo910Q/ZnBu0K6NvKAUdEzLxczer8FkAyisMMfQg8JD
pdPM20in1HLzEEKK3rNUNq4cxkBShoie4kLCxO9pvBAO6+LVsYsf7LGnKDLV7AKRt6HIg7ysYqSM
5JViIfdTQGAj3fBDHhcyaEDwiQtC3wCE9UliK5fE4aqn8PgKbidMn1PCVPRnPM0Uv7r29ZGBXgn9
+O92oZk02oU4aIXmTb1Ir6AYvuPSp+fmbEzT5Tctfurjb2pal5SLXzsQg6WVazufQznqaFUwDxew
9BDAmSr0A/bhzwT8dkJuT498PXjC7btptyF2/6Uq2fGiQ0DguWgmAa/1wdt52Vbg8TSaSz2quqaP
DOuNpm9esgreJzcKbP9bcx2AFE+cGGxstwl7UAIx5pADFh1Rp++yrQ/V4AwxgMRsU8iu+6Qir7Ss
Elbd+OhBX19wFNnSm8O8mbo1KMmKX1mctaXe4e+eSYgfJhs/oImns5qckPmPryeO/4XdZHSSxBVE
DvgHpq6NfRNCxhDYqQ7DXfT1h09L6IKqRmUAZoVg4w5prEavOg+QcvwtsXHidFAj53PpTpagNNVU
zW/wQ/tXrqmTu5FBbwj+Ero+atPo/VNlg+NDlB+4nu2ZhrkCHp3LeiaklA4duE8+XeP/U0CumGVq
7WwvDHGcW7U+jjZOzH2YhcD9yaC2Flf5Cp2qQ46CKQ2qR69Moq2sBM9O4bgZXLw2zQ08/HM2KYDM
kfyTNk14zcxARXy6+VcYOmNZDIQiFQ4OqfoaCx+meHj9xVnmVJs2uD5KcH1Q76lANFmZtwXRb6d8
f3omiYCP2urhgErJBMXWGHFGepcCSqW/ChntIKjJpuJt3GylicFkXXp7Wn6UmX2q4YEfPrZMODVV
woq75Nyk2KuDNBHR3hgIFqPgmgw2ScTXDFfYot6QS+w82uEBjtmdvxZA1iP3SnDlQvtxESbx5UjW
ddJOg1h80iI+EZ6SyO4RTJSLneb+Lif8jZj79THgZLeE6cw0SKKIkpN4lsMamOs+871zESiXQlC3
a5irLRVnPJyCy1QjgNM1ww0TvG36oibUeXzbgGMoJHo83zbHtE1AXZVyJ5dWGFqe3e1Ykn4n0FoS
jxRd9pr8Nb6YHcMFo2+pqPev9QJlYzFLcdRC9GSUvbG13rIDWkgtKMKTMLD36FJPpTJVTeJ5ipBP
QTrn/ez8F+dWge4JRyYyGVgPePpWmsd6qsYrrGrLIQNOr3FAM86yATRlFJMptH2Myin3JVWXw40X
O6sR+ucSx1nIdKuqZVXioIXlzVyiXLdEdAXfmFDeHow+co+5T5hrcg/6hjq2+cmwAX0QckCUV6yn
jxxaiymRqZl2rHnSQ7ku2fUVkoYgt4JUntSdSNOHu6HybKnWBKM4JN4G27k0TO84M9l7UXO1/m1f
BH7T4Vo9+7r364PiDsqvedxphKhASwDohSg1xPhYMikiZ9GpWpX/L9LU0kSajvjDkgHTB8wzk6oL
cBcv5LujXCs4khbLAj/fhavN1HJceT9f4RhKoE+w9y0Fef/fHGjmCfvnusRnsXe0Lnx+IHKwZ2bv
AJYJf4yEiMN94R/Qwd/UgNa/xUCpuoq2Jl5+B5Ouz6WQaHhtdacos633XcIYZzcw1aXkbNzN+AzS
fgveiB/OG2mta6JbPOtOZsBpvn3op4N6nZMcw2f32MRWI+OwVkh9IR4bMxfsrMN+8iNGjSWIsqZc
cdFBW9540vNg2oAY2iY/QIiiFAk+2DCrsyMDREeMzUn69+JGkJn2xUKZf5fNNM/5C9cuRYjqrbdH
EWi4v7JQNSAr7kY8Z8tGfI7gioihXT4ZfxAsqeFatrVTNCcJSsz/eznJoaVOXL3VMOvOsI0yWtQ0
sXMrMPgert4xD3p7cS2o+DUyJKpRB+NXOixSCWbXPMJlmABEJHbJMf5rsV7dMvvtAq0BqXV3gpNF
xf4nUbfwTpeYFbB9jUhOShtLlWF9nSudwKuatrH7JfjGaDTWvQMZhlwOrQO2HxSKe6FeXnmFwMsX
C1awN5WdcDjLp7Qi97yBopUffIooFHC/PXKH3Hi1ZrDZJ0/pEhpjAwsmVLVxVOVTfCJ9/do6x2J1
bYa8YHqC4YeIQ6poZsH2FNKffShHX1I45HqfpxZecQAU+zxLK/sQ6aAij8BC5l+s5KKGQOcbvbhC
W2GtKs4f5lKey2742EIAhGHB49J67Kihj50o0WPL/N2g2gAGQSa0MGIxS9gA739wg3i+R6RGNZ+D
H3Zkkgcn6ZwhJCrVUavxMBiM1Ll/Y4G7ebn1ky4GOyaPK7UUnk9FlRi0C5RcXDjPpKys3GBsmNdd
VwU12tBD9rYCrMlXDAyWnyNaYriGuDBWNleQByNVMe0i9qsz0DDR0sY0cP2yd0I0sLAdI5X0/7Qw
DAH2IX/S+YPIZlElefsJiQa+9T3uRxFoJaUk9dP2PR20IWNkjGaGWtspAPdlsYK/cOgwRNGGy9z3
mpinG/6ZR+FtZm4h5w/jzvcwx2DrarItyKvu0bvPtWU4EsJdQUPHvEx52TSC8T0+1YnfXInVlIcg
zvYZBZT+A0Vq/gXXKjhhXm+qx6XhVdJrBcyny8lHVWaLh8zqVIEK8u0qHfudN2oivKqAZDy7Y+cH
FObq2AT2xlempql3cxA618SoFGD8nITv9KfVFxXXdotPELJnnwK0/xHc4Zbgrx7Qz/I4qV7qjZkB
67eV9tFCjnF6mjhHEKvazM0xQGnCKWq2ZMoBpQMRCxY0oelnUphO7bcAzaJv84W2+DwRdbduSn0d
TT4gwEy7C9D3sJbJLGMKpc/XHdfCcFBAOUGcPzLdFJBW3KzLM+t8BTphs1Cg9Xwshv9PfXNaAwYI
mxReVmdCvCq1muBUSIGeV2h5vLyeGhjONPAaxd+8xppAoLwB5XyE2igZvW/sYvty/3G64MwZeDNU
7mj0V8qpTRnuF6i5O+MtG5SwvOMXxMhXBsS0s4mlYx3yAaL5X3oDInSQcvl44+giHA2+eThXDJA6
p433f1bcjhmLG/yRkMFKGoTTNZehDldhLHp/fCBDL5RSOykVtkv+Tpb5P64BVF6vVsRF9Dpi4U2f
vfH0HC7RpRguKLYnF7SJlZyhBGMyVPC0oPS40NWJvm/x6mh5HY1nNYMOpor87iJh3GHYt2WFpsN8
bg0be1G6wUArxF9xnwAx8ZzAb1Xec9u9iio5tvBIQf+QlrvrIL1lMN1M1bzjroUbvykfuvHW4LOy
871UvrT6Ptou1VRn50eMW/H2RPyWzSwMYajYdEVsvQoXr82gE/3a0Sf0kS2uYt50FuFc9lIfY/7V
bbf8L0/ahYOyxcFbOTdnLCeoeqHr8dPRAuog8Dn7gB565EjVIMMlvF5uAnQ1NEepwOE591benA8U
IA36ot/nwiPidcD09PdTPwHP1nROwJONL0Rp3IOKN/Hj3QSd6FiK9OExbMAAKiZLRYRNRE1K9Ct0
OtqLxM+zXbjB2mkpCk0O9c2PnKFUGw19VR/aUgkX46t0xM7uV6ppGTQOzlswPogYjQBsENgoCn2E
ZLk7+PVrRJPC6tcKyza1Osp3DkNW/XDMHfSrcDoBELuJd0x14Z8mfdBPgUNtmveqM9AQbUy0OcTs
jTm+FQHv7faqcaOUvqL5Eops7pBfVspytoy0a2hL8wwbdcUdAa4pDq0LAnmuFhbhEIJ5soHDePU8
hULgt0lVmeu1oGIXiAXczxEAIVL2tO/v5YMXFlOAQeJSu6LzljZxdSCQG16HPF/uB++nmATFRond
9cLrFmouRXW4TDzCR7wnmSGHzsLtvJC3SX/nCAusdWqqXAh/khMpfnhwjC5CgRYswkvi3UHDz0sU
9dyJ2W1mBdGHUri8SfJx3Aj9CQh0NzdaccSwZaLIkkIngWcsV4lof0G0XCuVfJ47fdXETcmL+HlK
f97wfw/rMLWzVsWl6RjZlECFlgWvKyCv1xUgaAhEotUz81NRWZRnkprr55iX4xYfO/sQJDSUQwcW
+88smm2Y3pK4ScE6fccRykWQDKjfQigZTcPiogeOHCuPrbTgDACjHPqizsKoJkTnWlf3AdNZ3f67
6AYrAkqCAUQFD6XImb4AVdU9mOUwb35aRdLiTtviPcWBu+BrfmVBNCsP0xqgnykctxYsvXO11SXQ
gKgMhUGX4qLexfkrcREeU6yqoIRxOiJnLrXevA3cLu7vbFSUT9XzAmVDri6eZFpd3cEAk0SJbtSn
bTavze277Rjq6Tm8pxlK90/kJcu838EZy+zVhrydS68FrwHrtBXqNSgbAwOUtDM33V7u9EIKx9CE
LsB5sxtngkQS9SVIzNxORmtlL/72/Oep2wCWow6V47zy0Ug3KALNiJZxfwZ6tvYFl464PsFcFa9n
77+21VpoFPbB3cRICCGS9NgYkwlged6QBVw6k76QTociV8ZWXhmushf5g5M9DTTeDIef5auk4fLr
EltU9nMs6l4IwHdhe3jVqdXOfulAGsI2frLMfslviBRpacvDNAq7E32/PBYasCSn88QNh6wG4XZB
QgtckaT3o7FnaaV5pjwhXxxxacUmow//2tvWJnOfADWC7kNrqnYyi9OBuVvtQS19bEnYffHwINwC
NoK08V1RceeGRG6jzlXe99ENaGChDofHNXnL3h69H4lWSEth9gXjs5/dcdfR4sdgK0ClNZ/PPcdY
O54ZhzlDWq9Md7RbQVhLvkVZPqmlVlksHbQzjT5WIEHqShn+eputVpi/SZ8n6P6bUSg/cvItDXvQ
eQOMSLgSjmee9pJNLoucUoM+7n+CQkq+/2bzJn3Ro567Mq/eA1voNxM4EIwA4GiZAck8gkrmpJzz
A2eesJ4D28JJKLKdG6jD7WEi6/0h6FfAoALks7vkUofuA8QHmXf6ZPDtbt/mpDMyogOoVtM4fMyI
7B0g+o/C6r/RNU3WRU5EY6fE2tsQWDaakhp7gQAHiWDbl0X+gY9EbAY/YWHu0XfHTPUeH89fW3oC
+ET1Z1vr7CPf0PAknW5wT9ZYt/xvtJyxp2kWLBLSj+jkUy5opx8RkDI1Bi07REfDoBOz9qvljpn6
iqYXzXtAGS/tXKSPfcW3t/JD2xoqsWsCQR2xbLl+gcpl8IK3Wh88pdflkNV/Rf8RzHT1Elvb+L74
ck4wBmwpUJ0bmkfVhzTSP1W0E/0CuUbF9aaMCBlDgJdQkAOS7DRKWUo1Z9PjMt0CQufFinWlK1zG
bQsME5FDbenms1RTnefUokEskdTBKF58WjXbbSl4jZBkxnpwGfH8ixOviN1JEumworNuHLLs826L
vH2jyy6kUiyvy8d3rwWZDDRCIlGrnNW+SB7E+yHQr2iddxqfNtXViWBKue8Kyzxo7CwO5JChuAYN
CfTJgg2/v0IlDHeXHSI+19MFlbUdOEzqEr4O7WeOjmoZMdlymUFoRykGVls2A5SIq+iMe9jk/L4C
Brc8i1AHgaNl4+VgCDwLEAysmJ56HBU37B599diXwiSjoFIU00LquZyCXfDX59JL2YvbcLfqVPEA
0oYr45pUfBUvw7L/aIDPKG5KCjXNIVFYWK4VhCScYlp8YJdqrjA7A6fXMyUCzpw76Y5z4pJT8icp
ZSuLpqokqglH/HqOMoWPyD0eQ2R5q4DmimjdcX3KvXrWKYCToEBHnvzdxMShDiOboLz003IMuoRR
eOB2OdUCetMTG1Lm3nPf1XnDlwcZSII5Avkfp0x8twLvRVMHV0N2LyEEuORlTTMxzAlIeNFFyahN
nQ8YF1y8H9hPjO1ZPxrxwx0fYK4TpeF0r+hz5WZn40PUH8cwiqaZYAD+BAlFWUWO2uZh93aG0YcR
CypXtr8hEkNoW/8RewsrEs9ip/113t64gqCbBgwQJCSN6eCVQaMBy+Xm5o1gYKKE1IhmSshMIONF
mNNmfQ5D0xuvz07M2m4gthh9atbtXDxJo3u4PpO0zJ3NUiFcGJnGgQWGBocqzZX7tN9Lc8LkEu2I
DNTzSBLYdoqwfR0LBFkZYH68lE+vR5X1HXtwr5bmGKJcC25UizS0shcrMVUN9Dr76v+sK+XhYyEx
12ROrJ1ooEgQse+iDEmmWQTyiNCNQM4YWKhGSO4ruMioN6+zIWYoTrOHLR9a7flkpCT+ymEsS8Cm
xVVLEhxTDBtSzQZVjo+IvCG+H1+hJ0k7Mb3QneStMjkapNQ0bxQX62qAz+nNTJvKbgb25euBOQlK
SuYaTa39DlBvjqygUPRFI57Uin/1aTBvTTMDIuR3PU8UQK/hG4oRIKCSk8B5u4Q9KuPY1lxPYGR0
4t+HNNFD7RojEMHng5/AyRyFjiwS0nBsyn7TrrXzn9U3FapvTFPA7nSXGr3Mtn2ddXaV2Z0pMblI
vMfTUuwxs3+l8RqeLZPGFX+uw42knoOtX3OG8n10nVoqsBMnAKTzic0mIYg22HBG/L2UVwwc1OCx
WwFdBG/aG3kXs15/0d9mmMjanygqwtgxz5s/QWXZNIfAB5ZPHKegb7UT/JmTRGeebtOLmiSIvTS2
iaG4MNuzcEAahqFjwqwe63oROMEWl4X0bOnuO346CZAv2EgsPCW4SQqjnDkbUAhXqryGlugeeNLR
6UBak3G0x+ZsCUxOESuLCTBo7ijPeasqJzwjgZZn5B4XY71ObJDMMFdDgigKpK4SME4cW336StJN
voltVqVOTwt1zXZtLUEir2AkHNghaZfGrQqX38qTY/6XO33Fr4a5bnPGDcXBtViXaI54wkhc431h
Ryl0A9u7d7o6qfUCkXzaBY1Hwq+5P9kFs/Yn9yLZl6v+SHHVDGGehWL1drsf1IiOuK4uRHgjatDX
IR6dm60Pi3xatIGgzw+D+8b4aReeXf8ZIpBEvNKf97D2slLFRl2LyjhG+xykDhOb/sLymyyBPvyG
KVPd7SpeB4QKeQLOQ19jwlm84WQTtvWKFGExV18ZEitcm5yAVKTvbf1KRU0/5CJQIftIAcXruGTd
2UB18twh0kFxaajZ0rGoyUxvW2MDneuWulcnUcmbPsPQZcpN9EhXYQLp6ApafvmaXZ8H1nECYEy7
4OgJlnx6eQcneh4lJrpcQgI0STQxy9eJ7kR0bBnG1jaT8cBV5FjCYNqz5GMMsDMbC7P66LRC/kQu
GdehyEOCvU8PxgZu69jlQq0eeEzVLznYuDNd3I7RJASIZZ5V69Wgx3ao/1yneQupvuHQ6PcmFJi7
QnZLEStdqyrc2PJQRPeyOU/E9YAm4qrum0b4UEBaRuljxD8r902xz15IWyo89FUe3A1bW4Ez7aKQ
TmSWZYQlLQEekJmhALvYPX6iPTtNsLkUF0qIca6ladiBgV9OwMEdrtPlajxG9eYZeR3eV7P/TSpz
sfui0hpdA5Vq9HJxKRFA7UMmRs90D4yEN9KpchDxZeCIUlnpb5gb0DisYb2Wk4LCDth4D/v63ks0
7eflaMa1vnpB0LsdH0laPGTf6we8GA15C5gT/lRyRDBn1tBVNKyPTx0Bwl+Oh6MQEoCqZRAbBrHa
tBERDqSxG95QEA4wlK5gPmc0hhu/MTgxaiDFLyz7cCTRBQ5rWuGqVg59vavvm7nNsIQ3sQ9fASbw
D4Mry6dSxhYACKKIBISwQUHdfnzJFMXdXaB4HfOWe9U8mNPIghZLOZb4KuPbHWRzffB7DDP//U9w
E4oA1+C33wWx2208e2yPep1V7FB7KacQ1h7SC18V/6gzJ1PToakuRxF85bB4YikOG5WEz31oESVl
90dRpdud7VHqLWNW97v0ND/Zsw8Cy6rNVwj3zoECDec8QQhZw2s/3Uoe01ShYllRHoAhfKkqyXsP
Tc7CPXv8Jh2WBGduYlRDUGW2vYTXQxemgXcIhr1bsvwUxR7qcJ1iNkUV5KKsdxer5L0Gm5+/C/n6
ot6KAOoaFmxn8R7oKWf0m8frvaO1srkNlfv6P3n2pWn5COjSfA5dPD2qY7pfUrBityKvknx6kxI4
bPbRqvlLAIFBwkrFx1cwMZDzhp9g2STi8lI4f7ya/7JkI/FznTLe1d9Jn748CxR/ROYQPfssFUdB
iA8wxrPy+qLScK8t/UGFw/9byxMaNYY9EdjqZN4b3vp8BEMA9KLhISRLkoWAa2WidXGgg2YUpfLJ
fYtvEhgwnsrSSNlGzRU99GOEmS7KkbVND6mSo+Ach2tef1JM48w7612VuAUGPBjaFvJJlPkogAGX
nZffFoXqPDJxGYKlF3ADQ5ujHgEIiKiqC3v6vw3hRkfuahfkCKqL7rmaAa7KKDv5dmWgQCJuEWto
AjWA6OdYn3NBmIfqpyfBtE5hFzF4swVgLrB9L2180GqaeYcQdhkrbOZl4jbsDwyvF4C2kMl49HJ6
gsCUa5egKUVNyZe2J8n57I0kUMcOKw2Xe73+T33fr4niP7h8U8+e3qlVhTfhQ0fvEDF8/E3Tajju
tKEi0+gl0QoVB7jTr66PT8qqxJDup8YWM118hv6oKn9WrjTdehJD6G/b2lueNwmhv+S0z5jPO5mv
aIrupu4hGXbul5m3HMRyBBV51I2uvSM5T0KNzSIitDYHpOGbLHcWpox7N8FLlwcXW2ubdOo8gt3j
TWxLVmloZlaOyACqIWqzfjVPpEbhkHyNxz/k2EfFRa8Rp1/eMfBSGzvRK1pc4HnaYGaSWapWksKS
vYlTdS53RiWYSCYVTja0zMTv5EgE7abnBWAfQxGxbz4Fl55r0qtBRpgzKcCbGcvVZ+RXXD19vzAV
GunCqgoNdY2lUBBOJZJ58Koc6UdklYSdMLzHDPxX+DPy7hC7njv5gx2zuEYYD83IAyjzDAix9K6/
ebM3pua0SpSv19GUXVsbncGsUxZqQJiqo0EX5YKvZ+MaBLOlRcCgB5Y/WMtztgeyRkNuEl9WZ4fM
8D2fDRr8m5IcU6kVnxdF31YoyS4s1otVbNbYK9u2J2HJ+k7yw7qxk+xy4x8Sq7l3PeoXIR4DxYCw
RxG7WoxUFLDvgiACkLNKoaBdgUWv6NAq4Iix2mW4ksoxRGmSiG/qfpgJQR5a2F1Dq/tpHF5yPeE4
qgN/iwom52zQWYt9JtRQenl7+dWWJuCbmsUr4z7iT8xJbXSEwNSJG5Tqp4ozOyQUKNSeB+SwY3yg
5lo9XjU/C+X86I40zO/Miy3TTQZUb5HQc8Ol+4I5dzRRFTC+LO9h+/cNa2l0bXXS+4zjZykFMeeI
P5Ym9fNy2mMJePKWDlHqmAtmUUeFhaY81lHTZPupdoaVySKl1964tFCAC5MRwp/BOxDm5W+q5+Mm
Ha4NzS9Qek5bvhN0hAbaRo1pMCkGkhySHsGrtW4m3SBsIsUWT9Qkef5Pp7L31LTQxIx5xfzaqhc6
8wH5Yiyk7ZmKzZne+z7WFMtUZ3gi/fysvCewGHVXS0xFqsDV2VUUmK2AXgY5PMZbTq/whuxe8vfp
Oz+LH9nuDBOewSnLoHDfavv2J8ZkLkUXRtWDVQHX+B81n+eXmKQSxWMTA+QUIhDVYfxQ5b2joVKu
T5R7SGDtqM51Q4wwLHjAUO7/s9oGtmlWp041u9BF2w7czWk5CcuSeVM9wTnZHexWNgn6YU50eyfS
kCkfhFPtSNv6MMpApKn7agHf1m9+cQZvBYhNgi8oCloa6gdNN7N2DrR0tCflCQnCMwn6UfdWfsQ=

`pragma protect end_protected
endmodule