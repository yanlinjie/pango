version https://git-lfs.github.com/spec/v1
oid sha256:79050533fe3c031089b4a3342fb697a6f6c48c319ae2f42851f7d7c827ccabeb
size 15784
