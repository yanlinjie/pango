version https://git-lfs.github.com/spec/v1
oid sha256:e75ccd0b9fee74c7f7db814116421a0ba3183d60c2564c46712308ad782287d5
size 1500
