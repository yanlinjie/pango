///////////////////////////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//the trig_unit module, it get the match information
//
//
// Modification history
//change rst intitial value from parameter,2020/06/01
//----------------------------------------------------------------------

module ips_dbc_trig_unit_v1_3
#(
  parameter  NEW_JTAG_IF               = 1,
  parameter  MU_PIPELINE               = 0,	    //0~4, EXPERIMENTAL
  parameter  MU_TYPE                   = 1,	    //0~5, basic/basic+edge/extended/extended+edge/range/range+edge
  parameter  MU_WIDTH                  = 8,	    //1~256
  parameter  MU_CNT                    = 0,	    //0~32, 0=Disable
  parameter  SIGNAL_MSB                = 1,	    //= MU_TYPE[0]==0 ? MU_WIDTH-(MU_CNT==0) : MU_WIDTH*2-(MU_CNT==0);    
  parameter  MU_CHAIN_BIT              = 25,	  //{mu_function,mu_bit0,mu_bit1...mu_bit255,mu_cnt_mode,mu_cnt_value}
  parameter [804:0] INIT_MU_CONFIG_SRC = 0   //the initial trig unit config which the jtag still not available
 )
(
  input                         h_rstn      ,
  input [1:0]                   clk_conf_trig ,
  input [1:0]                   rst_conf_trig ,
  input                         conf_sel      ,
  input                         conf_tdi      ,
  input                         shift_i,
  input [SIGNAL_MSB:0]          signal_combine,
  output                        match,
  input                         trig_mu_neg,
  input                         conf_rden,
  input [4:0]                   conf_id,
  input                         conf_sel_rd,
  output                        conf_rdlast,
  output                        conf_rdata,
  output reg                    test_reg0           
);  	
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity", key_keyname="SYNP15_1", key_method="rsa"
`pragma protect key_block
dsISU+cd8DZEMWwAWyg5LXdnfAspzG9KoiHma4yv84bFJH0azt/N1Nm5q2TAsrcIvcZJGITqckuk
tLn96KYJW6lOOxOb6IDC8lQpB0ZT8tvabBMfwSf4I0kRVnUSDAkI4EDklJnYoKkqxEYZlxQ1xhL7
8Lr0oKC3eaQrwMcAn35cU9R/Sp3N3yzT2dazvXYQHnC+HoJz2yPnTqBiTzZ+Q+aJz0XM7qYCz/Lf
7R8xy3a5gppz7mUvkIWXpmj7sCel7A/ZY8GLGMOXzY4095GH7/HUL0jTJaTwXihbcJl2GTYp2jvj
Fa02Dm6jgq+XdsYKm18UU8nUq7nm687ELxy/aA==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Pango Microsystems", key_keyname="PANGO_V1.1", key_method="rsa"
`pragma protect key_block
IpU0Fl1MepyieHFXhU12n3O4vG5kx/FFhre3pxv54Y2UOpX/obDh75VDdu32Bca9ltQnV5psolio
+VXh4owkV+829ufCdTiAfwjIygqqjEtMwM2EEOuxJXAgt0od3Tx6QlZEXwTagYB/l+Xv78o1a91Z
a1bwe0Wg/VEDp6VRekgYgNYhomnkg4/arVl5uVy5TO8HcHW/w1I22E5WF+9XHlzb1Qg5DGuj9aaS
oZCcaXCfx8PLH4opldZ51ADLKzo+0qlsF0VQgAE4s69WwE6mqI4eO0kVIVvFIWCPoIj3T2FVS1Vx
/0IxXagu/l1JSMVngn2lTANLIh6W8MxjlQoIJg==

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=18464)
`pragma protect data_block
LBKmbQdbeaLM13bWyn0VfXo5rNswDC98fhhG4dOvX5iOZmrQkByfGyOoE+cIcaYAtsP0GWL56jUk
JhwSid1Ed5A9kzdoGo180BgXibIYFPsLapUcaNhLYOs8+eIy5dd4jq1Tr5oEUOsirjvz2rq1DI6Y
IEbBcLcF34AsdsyWWJyyYPf7U2015lzY0GKaMOX3JGnJvGKdXvGvizEZeN5W3hyrszI9YcTtfqoF
NzmSI+co32J6hE2hhKwyCuxr6zAacLoELGhW+u0CQjnO7/0f0L8G++OSX/rWAcHOuMavc+FPSMm4
3apbvd9NnOz2kL5VHNUcqsod2swIDZn4k+2rzya6LnuBaoMHhxrs0RshlT8IdbJixNixQSLNEGvb
bq4vjtyJkvcrNu7+MjKKpW9NalMH4uj0Mw/j6v5REqrz0HPw7qJhaTuCf+ZI8pwAfxOyNnLbHMSv
vMVI58+saBS/zXYX1bu7b9lTr3/HTr1kT7z3Ddu8sgNpYXc7tf+p5XR67UGhFW13AgdIBHlAvefA
MAttFr7UxObY/PkixwXJLWovAC/LkvOldvjYYfehY4V6zjvXCXqiLHea68bh/QLCSEFmCPXbTffA
RCtuEGaoPLEez6H1a8ocLKUUVGUwu1CR5msZIcTboxqPs+N2oscCiQokOwDXw7AAGRqR0nvIglcv
IUZg01o9C1nhoIMAe3Jvs0BF+l88eJdfb0MbaTHi7HpMan/oDtS7liR15WHmil7Bs1P3rV9+QEEB
bBDt3CVMQlAOfwnhTUKbkjFxgC+tXy/rKcnRdZehSD5dEwI38GpvErwIKdc+xjrKRaDrjudBgCMk
i8O8JQEo9bdPIQ/3SflX9huQbZfpWqSII4EZml/IeNYFP0Pft3KGrRvyhkz/UK8bEOL05TVeLD77
mF3IvywYCXTG+r7D3ILWkCk6M8N9d28g+3rkLmW2DW+ZC4zmicbA9THFG3aSudUka7nqaobp9ivj
K5jI6FGPAvVXF1wfNqF4TFTnoMKRi+CspWi/0r3BKwN4AevNS3f489dAW7zblrizrZGik5BUDfrJ
swLV+aCzLkNqWA5pL6onUwSpUPvClLhAU4pItNz4uhHN0Z2KV7yiwZHLBPai/8MK+CZh7KcsncLM
7NzVn8ykznI4AKTEZ1ogVKoV93Q4maHQ3ABQT8C9BhaQomJI4iyle4wzKh9nWu4ii79vPX5jk3yj
h7dqyMRfF2CQK1BcrtQ7i98gapnlzuBzGzQoQ8nkUcK7DPbyJgNnnx5hz8UA93TyhwB03cB4nlEr
SCJrgqmySwk0bdqcQbRZxF05FgpQQpsxSuMF948T/R06562sG/07+9BbEzGfkxHCKlVYUPiboelp
Ja7cTgumodUBvTKqZRVs2xZUNL+gpbOozn0RCKnfj+sqhzv9l9y80hf4RhdyFjiswr6M7IIg4Dfz
sxGxn26MnaLZEKN23/LfxkeyusyqwOgGkShngAZvY+eXUwxI4G5L+z3+EwUCyIZ30d/od07incQH
RvqAEchCmtbJElfhuS3HTxQOoWmUwCvc3GsmLHq5ecGryFUpbgFdkWCmPmIdSjqSZU0wYgPbYtJs
LsNApuUWpOB/L+FGx5zJbAqS1iFLOXf6JXfn4zWvdjduVVnaQ8y8P5VfL2KudHPj3USUU5kxEG7N
NbcXRpESZxjlg5vbStNuRgyYFBVgphnKAH3dwRhzgtNTqwqhzkokYtD5g5yukqsVSahGejhwqKco
VOhj/QXlg6i0ewfpOQvp2CZcaaIFerdReJgnqLNxLh8Ekel1JhhHVWYvtFdxJZXgGfx+la3Yg44J
vJmzfwSjxz1IA6AWyFft3Fv6Co06ItqtuAcAjlDZracbZqXoOlciA9eTuqFTEGHg19ywGCDyvXsY
xVjm9OmstkLWNxlYJDPZJAgf/8LfBaaLExymhsl3w2fZc8AtIPMlEVLnx0RC3Ym6/uFf5euTfuUI
WyeZG/4p4aclygW5X26riUwgyfk+zEJo26+beDASMjd7PcdSACevq2md2kX+t08ip2Vg1wJC7nQy
/T8OhOuMIKsE2Eb+aE/P0dXPnBEgOvYkKsAcM9XRdwrEe+JidPzfgcX1yWNWDIcsVriUJ0D0c5zI
UBhyYo0i2HUTHbdJ0w6dzO2gRak6czWbhntUF/6hoba3fWupuIRerJEtx8xwdRS1zvf5AaTKK/6W
LMXfWGCBH1jRjrqLzeIAWT0MU2i6byU1ADqmeSFUkj1OeW2aV08hTAfVvcXw39fHrce3qL77e/jo
fA0X1AxOJGfXkqKvnlOfAcwDfxUsmdyIEyWDzlf/8Z2sYxNcsvFX+nOlK7mJgYSPJqEtKkFnPvVj
o9M8gW8/yIz7OWWE7MOCC+jjCn1XTjebJ7l/STcaSXpF5XSuAEObgyZVgSryjrPoJBMvAQ122BWi
OMLN0VG9jJgREhl6+EmvV0gW9GxOiycXh8fcVX9kozvMpPCyPTEJkVHPrDmNBCXZrWAkmH+wyaNk
1OqFwCuuoSnq+MNKp0sxCt5q0jvnG1jcQDmxjYdRAPLEALQx0WfRuW9quYK5dkMOXqmvtC5SwUWM
mOJocL+pqkwtGUC2SYjAxXI7HicsT5qz23LOFO/I2Q7RkqV7iayOe1mkbZymaVMwdZEKsxW0aFEo
HM0pwnk5Z7HaJyGR587Tw9r/F92yntGop1lipiITtFmr2gke4RvK+ik5zDEk1mQfTC3Lec417Msw
7VZbGmCctvtR0FSIse0nAc2qokoWH8ngoSG8D1KyG/j5HRx+hEffEJ1oqsc2vXWKQp6dQD7qaSEj
TK6K60XEWVZjwhmo00N9wpWyAkRrLO1RMnNozfYfw4yrFT+cwdJ31xHP9mWQ+L9v+ie3CBdLcC8J
7/eolw7TuY+f88neEF0QuI0e+UmcjLXKO6p1qjdp0AikONJCKTvC9qQMugB5HWshsbxpr9Y9Cy4o
KhJAAleUqBsthCwL6VCjLCS2iwCt/lMnM+FTDV6vyCMkEjmTcF0kV6kk8oqXl8wRQ7f2ecAlFRdb
DAOrQpXDuHoUYNORe+SPwzHzJRvm9gImDYUXeWMKrMV4FshBh4WlHAoS91pau/WbiclzRA0pPNmQ
tsX39/GZl28yih47hjnzA8BO0NDogYaj1tcLdiidR1/GJjMWyeGK+toeoLFGOTyNjdAsuGIIXT+r
0io/HoZK2bSV7UxCz2y7I4kP54KluU87NvZe0cUU8RjhVODDd8eullpI2KHHsxkniFt+aAT6LdD4
3eHhyn/rfm9M3c5QOYkN2LPCRIpYTcqXQ+1NkBuDBc62hnZnImttVu1KAKRkqRW/joW57U4WYCUl
f7dpzenxy+mhVLy+eh+gO3OJpiwicT/SRaZF5vcfOPlDHA0qLiYvL4ugqNpIol0nwzdsf0yFL1J4
AfLtAWuBCwftK+rQ/gCFP1WRJJKeLTyontfITilLGdq+K7Fjhv3OjAzjOxW8YsF+wGdGAxHRibRb
V5RAYgYqBdrJ7sXTPZPGOttefLc4GIlXxcJs0rmoHcO0t99wSPiUSDD2gC5224FeQP1bxacbtIm3
dE0Fy29OW5lHNDWoeApEduXj/mpY6cYJF21FX81F24OqDH2pEfFx2sRjkq5RU+dKA64meJ2sfdD9
V2jaVIquQ+inlDXkwwONYS0USI3ldukToZruGDo2hMJehRAaHpY3TH0o0kFDI5DTPSDT2B658eer
Cy6waXWAXS+htsAaDQLeHx4KLLz+OBFqz59QM88HA68iLo4sZRsIYIuejt6Vvq85a7N/b6BCwnny
h+Yw2pa9fFPo1FMIicx6Y9Tz7cPvc+FaeQzJehjHfhAwUXsJya5raXD2WMPv1jqQmgZvCr98DeLK
HjZDg2xpEuu6KHV+/ybpDKEJPu0JDVMPgJ6MmLtPQ2x4nHPjVzAQZfyyhkoxPXlB/UJWwdfuCv1m
bM5BLiPIDIhPqkFq2hjSBLW5LsYTUlKe0IPXgt7miNCN75WIzEnAfU/4yVxXfeet7QVmBdiPA/Xi
HFB7SppZIZe1y3nMaCejFs3b0Jp8xp58GkufYvoTbHayIg2ndK9CNdR1MC9yM4WTS7anghasQ8Ou
xJXRndNY9AidCkHSkpFajbVxJhGhapMx0eH9ZlX0bhaXEYfgcPAA8kaPlh4or4LvI28lUeSZotv7
u5pZQw5tD8Tqm1cgcKPV8LwU3RmM34Z+1SRVSV/Do6uTzaGI4uf1sFmARL0F0vZ5Ae+FiN7aFy8t
MGK3bx7O9FDZ7Q2HS7RFEgoETIJJCp30264HNEEwCi8haud8wcD/cfNEz0OIYrkT2kr34J4467sL
DqlQE6ByxnUi6RG8ZUa0Gfb+hKpbJFHm60rjT3vv301eFY2QJkaLC1OqlpDHRk5LhENwMhPnenmC
sJELVR4TMEhifg+8l0/g6x6n8LLaMqKK87ZoccznDhkJ1Cmy7QkCegzz+m6ZKzIYXSGm5nBkfZuH
cp5m+AXAclqc980rebf6oZdPpKSmIuTMeD3LWIhMWAA5Ql92kSpTHPkCczshOdKFbHbq+T/OBRXe
nufqer1TZ54wkaPuNyZ3XeH7amTXRwdRzds0RjoA6lJJ80V7Z/OOt6PE3VNkab1Vca8aOY5QluOx
Jp9FMglW8PWfm8V5R2ZBTFwT23gbibl2q/mR5vfcds3GYDDXIzRILRdH3N8SUbEWvIpfrGnBumIn
KDEsTe++dbqRR1yj5RzsdDe/+c2SN8QPoVQixiIg3xiodCamiJndl4gs20JaKzRAcI01PY0Jg14h
Oysd83wE3/D9iNRsPbf7Pgcvj4g3QYJXfEycCXCCv34x5vMxvZsrO8DY18RGUwC8hqQaEIKZQ8s5
14tlUD0ts60hW116/r1SITLadTpYBoRdCyP819wFTImdj3350vowLh1fVxn/PFMdpanXDwt45NFu
aBlMHtfz+Pr44t7M9Y9MQwZsnY2629Hd2DhNkb2miuQNKbiEKt8oXXA60GYUKj+wX3137na7V8FO
5D/o2Je+m8oSok78PTlMkY/IMPl8HY3VKWDfJ8EbJvAo0H0GIdpLu7h+ixj7loif2bVTGUsZuG5Q
NpiXuzDwN0M2Ta9Z3ILMNPc/2e9jNZ0zltZxdd70pAMF7uTDSSqPkj3W0R1OBezY5xISDcrjiMBh
kStJKr+xqij1e4adANR9ulGwcAPQLh2ElDHN1VqmR480U9fn3ISXld42CyKCm2eafcS83T+ZdR1m
3Hy60gCVhsJMgBDmxVpEyfi7W5LZ9ol5Iop3IEIQny5XWn9fWxyGLjwzcpB45irzeECy392fM1up
orCzCiD4RAtEY+6Syn0NL/XqUjGTNrc1HLqP6jcdsjQuzx5jcSBoYt3PkYPk2l7eCg4zMSCpduCX
+35gszUjboetwgCJkGy0F6ep0b68mAnzRRqrHXG+ftb08rUhNuZXQkH0mL1Bdnp/lTMuOQGHIXvY
/OeV6faR3oktVwntELgNojRe03EakgBpEOZjJE3+Q+ibGrivdIk1/LnfMxaW91rxCx+upfJfMJBh
PbjPVkcYkKKO8flLqn88HjadAo3uRqSnpc+8I7mQ2waQgx0KWN6E7phk9FG98bOoguLXzWUD/dfd
IAIt4oGUcrGDGI5KZtKTroxLc4nIo9PUAnrZ5b9aJWNWAWjvV58JG/cQliRWg1nzx8IfXGsog7HT
4709dQFmTahvuLf79fMYO99j+9AH9nqbzLsAO8tR2Dm5PCQkXdz7CCyBq0cWZcpEf/rCTdSb6hKW
xv20GH0+jnxwe7jo6wRcdg76zY1kMaaQ0crTIs7kKNGoUv6kQWBjiWM++UrC0mJbxKrjmR6a3nee
pbEYKJLpIt8MXN8EXp2PSGTOwqb5S6DR5jL9iNG23ojbFoduye0+k4CPBTHaKVINppPF0BOK/Elx
rD3hUVjgEwTwk95uXuTlJ3kK6M49ESzlrkTB5gFPgK40kCoKHcjuyqd3EdEBNgw5Gs9hbqEIY/dH
6Vx9mqFFQkgsAj9vQx5WaepCzNbDHtZ9YcVzq/96f/ur+Vzeymp6KAGLagPTrhmsPupvzHjWA1QS
ua1iGValw8EfKW/UFITL5L42MV1aTCK0Kg3P1KUyEGCqQAcbxugPFul70DH2FdQVK/pZINRzkuC8
4fqqPIGrOotThtMNOQnc+ZeJvW/sBXT+6ZN6lU3jlDfEBhX0UECDv5148WVdqoaV8aid6ISqm20i
1raKW6xWxgc4wrTbGHQaqmTg/8jwqXQBGOFuQhmw+HUWk9hSnJ4qUICUqiwPbY+tH6+VuvVtAGeB
teP1lVUlCszCLTmjMT9VT+FncYeAIW8uMpk1JCWiNv56gAzDpU/LNUdZLIaibD/Qy00TcrNMNvbW
MG2T8OOiMalACYJZHiDfg4b/EWsVveMIAoSMqK7Z8lavi0jGB5HthL75cu7vtUJHjMV5f0km3CJf
boDbR5WxYT3ggclA3pYjliqfwef6wyqzPdiC2uo3uR5Nz+/18Wm4Ejfnyc1R8dUnjsHFf6J6HYQJ
o5+pRqZH3duhTY0Wvjv5N3IsC2+BYsxSmL6JPo75ysC10oFfazeGjsq/XyQd0z88W4qkXev7p3CW
gswVL9yVB2iokgtz/WiX2WLW5eWFxTxFuCX/MlYVOOg9qNDMK0A9bsMK5IdswhjOxokj9JVVM6aT
az61zgt/NoIvpzy9GX1uN5zPCEIsWDF+xUiborXawUK6tLRKs5EnNy7wc4Unv1dykcXSZAmipQD3
1lMk1MPOKwi4L5M5df+Q8Tqixc1702bZ0yfS/U2fVE9aNENWD6OehnzaYHH/kgBCGj0R7OaInp4L
gqMUTB1ntMhhVEEAYiVfWkYRkvChhAyZLVDwaGpeHsbVSFH9ekzotmz7ds8IZNK8wXtKfBvTrLY9
4YDgbns4cZzTcUrvNBA4rNeVa/qzH6bbTu0ySRw/YNVBEuY46YLM0Hu+7o9dH/TVp0iVcVUXv3BG
7ea0+519PL5fW9IEM64vvTg4kZ9YxBs+7FXeOiVRu7UHx1zgmgO8RFDmulOePZIFTdB/xwLVuDwm
nC/CbITm3AZ+gRgUfR4TDo6NkZqkbqR6v2LD6DL+RU2Kn332gWZehfsrSVm2O29oTMrHsfhgdVJR
a7ulu1jHGKWoBsLqpomri5Gizq2DT07eArIzJ7fpIflPdc0SdD9fpmVKyxoDwk3H7cm2Wd6vUGpt
hqLU6gbzKlTSPcuEScJ5n+uvTo7TcSBFvdw9jP+G3Oih216GN0YGzlERvKkO9gcaEUz7B4I2ieya
tWVa7oj4iHgayOkImRUuGRFlDKxOCDr9mOw0PtehuWbWMTPTRL1B6s1y50b3byx54uS4tapNnw4h
xHS5jHcpz+RhmUYQfIzFdiRCgc38PF4WXe17V7WcqjCQUEoQV9Fq4ZPJCKJRjQD2zhjrHUyexiup
B+57LDIzgDoApsUtyRbi1jU+i5gB65PWdvyHY/KLrlpjIYhbu4XE5rXmEkiNpORlZ3H57VM9pB6I
6t/wUER5PmEXZyrlJLegjOmzOW7Dk4uFniQUqv5gWRwnIWbOxzqh44rb35t2xU24C46cSxMkLcpx
Q1SmbSG6Nx9Jpo3khkWt8NePlPVj+PqQfa5EbgBGvvD1IBCxaGzjttj8g/YwBO9Lq2wTBnj/CFzi
JGqYWAf4UIFDgRb3dNARsofgU9k/8jy0x2giHfLVN/OLxHLV0NAZvT2Jcl4PlSM1YZv+suKcUeF8
6Fba5VTtGyLc8NG59wvc62z8a2YCuR1y4qqzAD/YSPNUHN4aIgNlHa8VD2YFiIkpndkZn1gI6I6l
SXAr+D3lfPwe/d65TEnCULJSm142w2AyKYNEEtm5XucEz8SnWSjLcc0uDxopoFJZaJRXJvq6rHyu
rHtgtS5BlS9zeBaSfB6JbKIM3proAO3Ab1u+Az0a18BFF8d++wRjrCxj6NNutSgmca+i0uzmairA
GorYOVbXjH4mEBL8pvYlBUlEbEohRj5hYRjhjDw/B7YfxeOtSUF/YAA+qy+JdUgPwBkJgDNIiBc9
FN0qatXUBj9DwomDRmiO0YaH9QsM+2Aj85rbaMcUTh53ECRa18RSF9qGJHfrElBLjyy63R3INXYE
JC5NndB82TDdO+qwhf0jwlgTVv8r3A4DqiaPS0MLz/wkEfG+J3o7kJLmQRO03vGM0WDwKpTM1Oli
ZXXA6lbTsBH2cIGfC7Ht8XiJY9jdTX5oEhn+t8aGk8ureKPfasaSQ9cF4cS87jWNAAS/M+OdIXcU
wvKL6ELybx1LJcelZcZVefhATPsvbsBouFqK7m1BVGZfdk3xYxnKv3ioNW/6BQVpuZP2jSsZywFj
KNjMs+rnoyigDS0zLfK1MsJCD7n4a3XJzPpo5Q/XD5Pt9ViYFP3HQsVwkyIreooViwINPdvktEhT
OyLKV+psPjEtH8749rzKqjWl8pPtEhV24JEnueXF1BmS10Lcwb37m73MbVT/pTg3N/UUWeWut7TQ
bBYVwcIi5Ca8zWNkV0it1bKRz5h1iCtnjTQb30M3wiOedg4c5FJvwxyLhNvE/aTv7SghZDfbEtSg
j0h/ulE6L15lcuVciP7olET+Zt6vwT4NAnNX9AZ59xTTwhReq5mMl0Cn7eIEqhHUjjQU4VHf3jvV
eR1F6xaI6p4uWR7hAaH3ayeKiqErwvWQzk1TxnkwTzoemcMiUNcmLpAuTdIfZ6dh3A0uS8aTdjDT
3Z1X1rC2QPu6E0hnkHf/UY6F/Ogrp3KWfaPMbtjS4ATaGH20jXbrCyaicAz7XeON+UGXLFhq25nq
tLwkZ9CLyiqTo2WMdYoTlMfsi9P7eAyVeGRq5KujVhzvOkWBmy+yzklO2zvi1WL8I/iN1SW2RzEZ
BDzHFD/YDep1R3aWpO02IeATjfWoEFgRzxOCwSLbNBmAonMRgKfovcLP21AgLxOBO4Bj5FnCyqiJ
O6mYv55B9auoICtt9nAH8RsELVkWCo7PmwmnCxLdcAQ7ejv+ZlMUYlY3TQXBHpLRpGn/NRvjAA9L
h2s/xXI+uL2wqaHBsLn09onKroV2HWIBzXcxfLDM9FXhvLytU3PREKpQVgbAg9OaM9+/bPC3iIWQ
Aln/Jp5ZxWGNRsZ6IVfN+rUQ2o4x7YmwS870aO+apORK9Ux/3zffD2ikn8/HQkIBqy8apGSnDaDd
rMJr4SoO/EPDoFk9o7ihfuvohiqPyBf3nVspukHtlZyay1om0QJlEVYW0I79//hA8YXgZDj4bB+P
lnvzYyeXOU6ywjUWBLJufI4xVT9aW8qbEkMAYBsYQHOZKpsi4HdvoYAp0f1bUCqRGEq9+INC1Lft
/4gTUI72jE2gaa0gd92840YMbaeZ7ius9wjbCKIl7g+ZFlc/NgEVa9OJWoflnmKURhshGs+UNmQl
iK5Hh2nDKOplvjFe6E7lidGWvbLTWZtQhkQtQ/PuOlX4KL+s/nWvU1kgrb4lXlgGoiIqlUdRRvgQ
qx5mIdAuvMEdpmsjMbyhRnqXZaHQLu1w9BRzgpudsp2k0MwXjG3t90QN+BNZCGWWGHGrppshs4ZB
EXvHSq2F9USYWqjlckbzRTcs9qVikwIK5U9ZML2IvfcvmB9BHG8XicgzX1NgXj9J3xBOSJ9BFyp7
moRH+7CDDwJp1+n1iZKb5pognkTnzo7oiSwQu9IAxu/vBc8kLhhG7LvdewkrtcdjRu+aZQxQy2Ep
oHDxRKJVC73geZX09Gz6Jjh9oLX8cMAUyH6b0TaVL+z4Jp5w/WShC3flf4fwmlMaxXYLXtelQNxJ
VXj1drVcYdCfhW2RHs/Z/2Ss9cSVUVxyTafnSVXj4w/d8qjqDgzt5/J4af4ZTy5SJMfvqfZP0itC
o1zlq4YK3lEzKBhoV7NF0j8qRved6sDdvvNhY0YaU5CaU4On0H9qi3OUzfOjYPnNlI3aGjPTLnqk
YDIriyguvmkcxWoEDY3X615cDYH/D6X0H0ETOVzABunEk4SphFsB1L4gmyY8hKK2k3VJ5gt9k05k
CzEomddUNsYLQhMFOLhL8dmmpfPvsWW7MfjzDbD0HzVQjx+oFZ1ROXVUlJqPh6GCNzschDcy+fOJ
zuxxAPR75uvsXEfhkJHlvfTF6WaFQsY6dr/3mDd8ZEthWdw1wtsfwIt3wDhQSsCm/1d+CVZfxGnk
cdxYzWca6rTBEJBpTqmQVrg4ib8TK9J20112osTzMaBhWH/qg/QIks6597ClQWWghpant58e4GXy
cL5l5o1vVo0nX94/RRR2z5yNd83XiXD7XhaeSBMTTdrWqFcFUjU/7PfSNS2i9EmqMM6i1b9f2/VW
cMW4y3nlRh8ikgpNuSNVwTDRWYARGvMUxbJkgj/i3fqkiu3WDTAhaYh6kAWOeELtpMGOEnYzmCwl
98KYtmlH5G0FJzytvVmDA5snjXkptfAKkpa/lypstmRwO5NJG/FbBgJr+2QhB2bOucxMis02kOoN
FD7o3GC+7u4NR/Fd8sRsmllpNOuYAI0CFwLCD5dSDEdefeooXljJeLcIPavTlQrKCh4W3QHQSSUb
rw/ijuKhzG6mZcMFY9FZhvoRZw9NDo95pfV+kJd+Y54uJ1mGzsJZkF45ouJes74PnNhYHm9UOFJ7
aJeHohj/DKV5C4JmGdjQtWDihUwXxjdT8t/TT+UNb8jKWIA8yXX4KT6fGUnhB41N0u9zgYwpZabH
RNOQhT1xwA4mf2dFErOJQ15jSrw5Ywv9O9OGNNY2vELXBgzqiz1i9Or/Ed4BKCUFh9qqGlJkVzoi
QtTNnlKOxbSzGSRmTHoCJuifbbTySHTSMgpgvr1NQt9EgJWoLdvEwxgeN3JdnPjo6KhCO506Fwvg
izlJA8i5o+kVh13b3K4JId+awGT8/awEewizAO4q9FQUF05XXQyTNxgvlAa8ZvtVJTBLVWSDjrc6
1m33g69ozecmYJLqDtRKjk18suEGN+W18NkYRkcxuK+SJCQ05zOE1IpclagmTYWLlJeJ+j8DtXKf
Mp8jZxoSwKVV3kAFYZ7mFjggr6+2PXwhrjdaoO4vNcG/QAY15jyTw/hQyYyXVmvkgh5/wB2P7GEN
WH+deHJFRHbLduWkaRWubY4CKxB5r1sFONQ3JmBKJrD8pYY4/xN5yZi31JD7yvcuh0iN6fEr+PbB
PpJmR/MuDz6dZ3HNiokRHhaGBHuZpQCPfFM1QwmvpuPj98AmEhXbZQHoKeAAstrTlsolRTGxxiKQ
sMpC2gRq06uHgWPTmVHAUyWn1DB3haLj9qcSkN+ww3WLwPMnrNcJsn9jQ1MpdmOomgTUazHNzAp+
ov2yR+xTGWbBGukS6XWcWD+nF0zrGTQpZxA+V8HvUAfsGbY65Px4PxNOro7wK5937NcTVpJw9kKU
gtEVVDaNFe/RoLHupoDDb++EC0fkzlkPmuJxVsfNIsIiN77qI3JO3A7Xhc1mllVmFlOpSMO8lt2t
LjRi0rm8urPVh9AojnD8JXelx1S/7lDNi7MNZUenp9rfKkXDMa2kiTt1pNCXc8d+tOeGA0xPa3HH
NOUwbwl18PNHgLztEQq1LLf0Klvj2cUCNMngsDgmDOXyHbZCedXeO7eL4W4E+hPUWze/X8XYYhZK
ctTIBt+GSssbCo2kobOU2dsEKhsiJio5bbmp09J0nyT4+VBZfq++uaskFAnnEAHM/abEu5ss0mei
1g9NJpofpTHlsz9dEjtRt2hk5SfIER0k9T7VCQJ5sRMBG63RxkMaV8Kzlq6OohZ7kvJvAkan8luR
a5iiBgX3e9WrzZuw3/qdtudIvunvv1pi86dPT3nRzgM7PFO220gEiogTnHUPjuVVuUUZ1cFp8D2R
bA5aE/unIZUWPu+K0iAsDHxltotGf8F+/0cAG/LouGhj8I2Vp4WbRLTURpYvKaqncbXrVmPCmpOI
RPSE8pcXdrjANaOLYn2RXRC5RC68rfq6xjRHc7PueokbPQKu0os3sZPHQ9QTR5YXAlVjontaVTzS
7mY64rqoTqx5BawkBMOflx0Jvv59rZdBbelKQGI+9ayJCnbkPNwNAjV41xZqV3RT/x4EHBDunDoB
VtufpSK67MZSqioFbBAii3V+iH75+FYXy2rSlv01hRBkBDNYLsybRt4utiebFntUoB36N3H2vRzQ
6cchFNEYEZsmQdV/5giUvFJi2hFFuK5r86Y//0FVNVkyJSX4UU2Jp35OhBflbtPpBCK8WT8R9Yfu
QWKZX6ruP38y9G5q85okDlAmAi7++1zoWUM7gE40K9uqZFlI5SN6pPEuAxQH86lIDsKEXXouk2I9
RTXcz7evuoKfWMFeTDR3kxMKi+kgTcYz/0TrA6/RzZogjaVhIKh7yjPPCV5Gq7RlznSq5G5/bsry
gu1MjC4Al2Ywt8+/fkLaV6DPZC1GDAopdzqYMcDsTF9dEyplK1OAIkTzbkB2x5dLw4FDsPKWZMOI
icOjWVVg+dvlB6XvjXPJCp7+kdKA1QL4OXPfIfOSUWOxnmpLZKvSLjSi8cWVw8LElBAt1ypFNaGI
UFTvYWaXmxwT+EZ7zagfcxASenPJ3JuqmlwZ7iQTpYUaQSUoXpGxfEo8/5XY3gWkxFh7rw+hg761
CMTDbA44FAP9i0HHoOqykgbfhIMQhp5cgesrQ1Y6ylQHxGIXsu7Z9FFT0zcGNIb4lqMl+X2uN/2r
Vww2fyggh0Xia6o8Wm/VsYXZobUYbtsOKexwF+XDmbaoTIgIvQfgb9BFyVOupPKvOl1ofazV/mG4
3SE37XWqiFDLXTIBt51eM0Q/Yfj8Z4khDWbNEegygBQiAnHm6VzsmZkJ3SukR6emldTdQQmfOEYS
loIEJc0ji0ByVdMPTe01oWvFcLQi/xxlmsJQ6I6TH3Qot0lfpsOBU9K++dZSFEblthAB7QAg8iOb
AX0c7gY2zbz/FrGVsSz/7fT62FoOsd8rIUil0zJaxqVTurD4ZAB208Tt5QV+O5eKdf1LP04g8soD
1ZfFDV7WorZ7QFVdmISgN5i3cx5HPHnnsCb8rZnQVyre+Szpfw1Py8fHO6lKADjRpWeUWayMJbOp
APAgew00O8LdVy80MGWPm/10Ud7cTnDGVIxiccTEz/zOiA5gJA/Ssu5NQQMZnGCVrdxmh4xz5E+a
QR94QumXItQ00pgiSjIes6xIp3KuKt3q6PT+RELofaJOIVudEoZfhBoSvw44SJuzWFdi2BfyEp3O
jra4s1m19zkJ4xDfAz0f2MiDFVIGYnKeSlqr0nNrOs87tiF5lFf0+p8EXysYelJr/PpJYU4nNqDM
HhigYD0V67QJAAlBD3sRn7Sqt2CN4hBrolyzc1GMJYmbZ6fu1t31Cbpaoe/56Ev25juvBKdR55Ul
lB8TwmjJ8KlKAgC/J2ZcGtJfbOSQGWdPuxcgBOVLy9HXnXdNidZXDLUJCs34ptSUO4kyR1KbN1E7
AD+nBkhl+42aF2gaJnehbrkOptFWogKI9yYYmqrkZkGOEz3C4ap3Sd/JFbqZ/GtN9o/OVzqblmP2
LwqImWTyWbd3j1pvSRLpfs7lmdDmVuyRgawheG3F5EtZ+tPnr5UqZBVGYJMW71X9n3N5frYUoI2i
nnAKPGwV7TbA14DTTrUfJK5WKoVN8kfc9+3C8FXq1thgxtSEXoiX+GCIGlDsJdHzQM35L4NTdi1A
ukpvNQN8QYWgPTsvLiRppDy2sH0MVHB8CpWhLL9eSLbV+OLkHRxNUt5pxnTQu5B37bpsTP2zSObD
NihFUZK7AFAz+SO2oKfUk80Aa5SoJIhtr+7ZLXzeyT7twAjLrLH3HVpQbRw5nHce+/rOlEOhrxIx
wVTrdRChvMvneIxvDmTwpkdDXm0ZIYYi+vIcJTwlqvZGImQHpGUgLgFurfjf4b+qx7/l7FuybEUb
lciucpS3KIHLCMeuJ5CmcAmMumjRKpkm692ypPUuihl9yuKJEBXiE9rg020hkDgS4GQbaUwSK2XR
yhKQ03oTGrTuUz6I3BVcJzi50aweH4e5mo1h9aN0XAJBddYmBlelccC0lD1VrXQIiCpfJ5oGGO6c
F97+xc4rPcr6gBOx3HPeaIOU3feel8KSi0ZkSG1LTLTrjK7sBzbUk0L4FM5yzbU/BellOVorgyEb
R60oRd8YKE4pzztCKkcEiiop1Io0FtqdDeae58LiR+gyVq8fklQQNrRJ5paJEE2HGTPn6wY7jN3d
abmBrXBlgIt7xij4HsuadwXkoOLCuWPGQr6THCXCOmjAQtlUKMQCkHCO7naiWKkX1IyYX82Me3PS
7971mv/eQYo97NrStLTjKrzcGAOwQmu+YH4zUvAmcte8GADm6+OEqaPS6S5M16o0sB74eGBFVi0y
YIWlReY7e7LPQROworf8EUrDvzBUoo9DSWod517GcbytoatTI+kdORZaNnuWXBz44veMjI905gUo
JyEKNXClc/1HEsaPkISiYbA9amf1d6rzEj9nsZRkcRdYTTyCeFxbZMDc7vu1RVq12ptQ87Sr9ioN
MTc0keapKfldl60QGXdzKB1Dv+l5WusreaO/3RqVnFV28icF089M7C1cxT7XjVVCgOBFGuP2dj+N
ccLbQDcg1CQV8GHaneGBQwwgYIe+ZM9bzbdrYEuGP688WbRLRnE8tG6BnZPqApcPZYf/mAmKIAzg
p4WuS1E0pUxN0Tq1279sKLIldUZWbDtOcbRY8rq7AUCcOJNloAEBU7I7cH5l6PcAKCj16Fkcmy4+
GJtqZC9TowfbW0XZTKq7ZCJqY2RvTOb+ORThkCKSEce21v3eV2Ii01tJkeZTYvWbhnXZeQ1SrcB9
nzDOH9/JRzsNNwE7OXTDaul7ZarzrZWEP9BZslnTOrzS5uztpRvfD0l9MI+9rP6eJtBkb+6TE8Ds
1unkDsu40gLUCZFramPS5g3V5V023f3PNVhQDzbgXg1tMJQdDHkTrxh/LTq1gnKXsViFdHPlxv/E
U6L+QnArt1oJPQFYJY5yoLnPmYBlvYlqT3Og/POGHutq3GCxTAicC84nFbO6O73BUjGqfC5eg9U8
FgWWmoiVohbH9sLGnlXhkR3t8V0mtQilkjgLxCBQfzsUe3jjWDLsy3YOxmQE0CTi+vh4lAVYEU+e
n0MCMxH+68cJ8/XV03wBwd0X0/Yhklx8oXUVGEUTemOxkKBA39Ch72hP36keHlMGJgjq5HEijkO0
e+dAPd6FB8ObdR6DzUbhXBnl3v+C6mruRCoiME1mLyLKyuNpxuXyTfdr+jV9et81Mo7Hvoj8b5Bz
3R9fKs85xCE5vmahEa0+VW8TRmpS1PDgY/Qrav4FKsXCruPEi+NdjRetV0JT293CSwN2dOctE61H
JqJ+iPqROjO7eBq3pg0Wlv1xpqQTBAqqdPRBi9JwNaOOUWg/LjwxtDNIVlh62MsINv/mmxLAb9xR
aoyAC7I3uvwChUpG53vHj2WqfY6+aIHyqO9k2oBhI4/W9VY55JHoaRCrkPUDWSPw49aRcysD6/IF
z1hwFRWJEKBUXN15ffK1MxVD9dTsPf0q1dTEiH57LPpqG/4iSPiDaVy/4dPyXlJ63f2+fKOzUPP8
GuCdM0+/uAIHExvmRoo++krJ8Yabzz1r2mMYi+wEaNQf64qkwghnSoG+7U/PBAFzrNvxSgJwLAnR
jHt7MiEwTMxpE9A4E6wfy2AvkZSiaRi2NGKej5eI0dGsS1Up5L1lVJwABCGhoph0oq18dBQGoBzv
O32w266sNI37/TZc/nWtXNkUQZYOGcZsAb1WU7Nk0st3Ugp8MXx4oM6tBvp2P5c0VaLs7rInlqqX
LPh2Q0XtAQKUMwgQKw36HKV1n0/lOdeL4H24lTRghj82g7EiLf/SLylS1Y1oabH1Yfb1Npd1+f7S
N2B+YzRIxuzl8+Ii8PxnSxHJ56DUuj7I9wPUTTUFMoKOCgsF3HF8iVnLXzCj1hN0uK0Pc4G39aaN
JbD8lTdgkYxlrIGLBv/28nR2WEloLms4477bp2RXtBFU9e101n3ADqdL5nK4gXrF1SUD+m9pqF8M
ExJPVYQCwpICVz3K3XLsaP/Izho9mHIA5NxskfkvZ+HLbUiwqOptdt/Woxzq4wsyZ86U6MHfR0SD
ONwVtq9V1exdrk64wXkwjDeZ29XsbI7g1icAVWxlQfUEo5vVHHFoJ+NeWztK9Rn1lmJz4tbdnmCC
atVD25ksmoSYqomkdKGQhEin/iXhNmwMn7RnD1dIh5+QRnCxiqBUBe2x/ODtd3rpbfhT+hUCpdFj
0KsJeYFx6tD4rKyc5Odh764GUHjXfydgaZpU3RUOwUPr+v2dcrY00g/L0Yeys9hFm7kfSiBbZpdd
q24VNQ/B31hd5T4shFRHf28dgFW8kO4N0i4k0KjVYGdtRE4AwoKqVTzKOjLFT/2oExUYZDcYBqcm
b8fWQB9ECf7bBj7d/osJdTOL/CQbtnkhq0NUJW/kDnwUNVAM4vAe7KaY0vYQnwlAumMltKvhpP77
+J9o1KHdvCnsoZDXNtbeICY5WXO6DYOBK/MbRUx+MukKjg1ZyPTZiAlT4RSO68BPYChC5g1cvtXQ
jF/YUIPG8jjgPEtjwqClymZG2rJepDouHJF1RLRQNNdHej2kCGy3p8abWhNXLV0DJ9ldHcqMrjMD
vKIQJghfdw/3BBphw2XjD54BCZj4VP4mY8EiTibvQUl9/hI17ZcRzs7426Zhk42c1BAnph+mIGrO
rjplHusG8iOYfEBbQYOJcTYKcGdCbdFgGnLjGlJXPxc1Ha+prHMi1RBoaWNhVIS8hEvsQ50IDr4X
0V6oinGX5FSrB/C4RjmJHTn/cBxMPnCxE314/zESyzfA9HGhhLzz5FQj37S4Bem7fYcC2jaBd7mg
JPqrHf5H61JRZHKxHu7ZZ/PPyLlqrVrCwNfSbmbRqLiGdD9D9kiKPa1U1ablqzc6ilQsUD+Awhzi
1AGvyptGLoIV5ObLhdeU72MsUgC/o/dOf/SxvPZBj2cG+WeOWnCmdFQBXm/HDBeFO3roNWpUTIWj
yMf4WA04CMkvXo9m2U+fw7nONLR9Mt9GGm5Z+tOw/X/9RjnJtHCmjZ6D8oqfy3vYZZ2sUDvojURL
AF4ON0PI5WYmpGGEt4L/A8jpmfvjCo9pMnyyY4SJLroaXYg+bnjKJ+2u3PMSLXmajC6b093gb2rz
pnFLlhqmlSAtC92YnQ2gHQEeOqKkS0MPmDczdAnjuvux/b5VZg6cmxhtQbci6OtQA0j5I/KQgu3K
KCwzDkLY9hSzdolSWk7kkhNMQ1Lhxg95CChx/MoZQmh6yIPGTrWZLeB8p5g3+suMjEXwadsDrvTx
QhRoQsKhBOk0aFj03vK/qtEqWF+ndns1FLDYJPOxpyg/5ZRsCXIYf8l+CPqVcY1OS+lg8yh5qPYu
gm/vi1TZPT+WzCytNt+SZXR5WiLox5KdehzkG97eCJNyPhpZ57K5tAfCpxRFmAQC52UKtUNfpnI4
xrnNO1j3h8RjvouzwRdEkFbSRF9jEI0UG2TDTM+uR4BrzadUp/ghG+jArHmaoDj4GSkR8ze6k1lU
Qjfg+zmCF5PUFfdGcs88q5aqhG+Q/G8nS2LtOIj+lYF9j6wpvlC/eK4dvLdyR4tLp3BfH8T/SHqA
XRYuXDkA+pEUKAvSu8d1Cp835kYv3aDwjkwrFLihTPP1FcZk0VGZL7srHz/tnv5gXiR+DpiDqSYX
/BeFbcFWush1vF8eKfgrWMY8fwqGUgakiIq3McKBe9dvSN2h2h2rdq0HQC7vs7Fg74EOWgfw1eDm
7IGDQucqYv9L3TiZBNhuxa8aicvJSojJp3GBcgduXm6rm7MlENQV7DJ6PcIm6CokadfAFQscza+5
b+ZEvRy4hb+hJ4Vh7L31SXeOtYKE+0f1s4gTAZsVoJuDsxhKc3l35fyiz+2VXkJePjEFCLuCykFt
SWj9F0BhdPU7nZbzNGyfPMlGi/EYuOyl0Fe/na6r8Y4RjDFKLh91IuRHRAJHr0Rl+0kUZk/KcMRg
EBx+gtAd2nimf68ivu9z3UojQ/T5uwMRVEQ2vSez2AQgsIMwqH6uAQIEndjtuuWzML2J3SnZJ8fd
zpFFHJ+LHsIQUqwAPIkM+8Zjg6FlNw6WSXEYS0p8V1yU8kV7obRYluPs8d0D3CM7jWuaP/kzlYwB
EHXQ9tk3CgW40g/cGRXYxFvezVxjzAIGFOyD63/LXXqHF52vigZwHeeGlyaZRoBDCDYVT+8IFoOv
FYcxya/eMzT0zkQdDcDFSuL1pj3kCaXzmyAwOsp8CPZAzOud8U3gjGP+Cojb/Tci+6cQUQO1pH5E
u8ePJS8i5sfWfDT2EG0e5j/pankKqkbYeyc5Hxj2VANv0F2Y1M6wwhAoAGztIAkUnFojui+JjFg+
bh7n33JH5GJXvl3Co7jkVGJELcNzsoAxVuVr6Cfj0lEHb60PV1qoNeju6zCrhEohCJQS/6kG+UTQ
4Yoz8FZNma7bSb4pFhdMl3q1zBoxrzIL0EStxPtei+uHwV3mB0zvaS2WaBErWr7DE4yK7LsHhsZJ
6X8z1pfc8JhYZqiZEEaQXdXhM4USjjlXzH8nOLEAbq1OY+DPRxCr5yUf3se5DlM2pCMY42SC74lL
f9YIZZjlj4ivP8v0D1eQH+FVIhL7+eLCXSQsEr8cox8RxoVWTGthtIUJCWw8CdhzcECI16RwA9bz
KD4RqSDLGmKBGFZXgraflvaP7soezHG9uD39YNDyl1hGQTaEpROS/re02cJqnky9FLUJnTVvSAlH
cIn90BJXMDLWAI3dO8W+LL7je4YXzJTcYf7Liud5E1aAWWMQ2ynO5DtzfW0GTQomLQbwJtTK4UMB
JDbujXou+q6IvosW+RMqVo+M0yMOu30+mM92gJXjIhwvmbKxW8k5Dig3Q/6UqRWoxsM0ZbIl+U+N
hFAG4y5/gmnJSa0vBXeLQn3RJQ3nRWx7iXLCgdpp88QAGnLluIpoe2yQkoeOWodq0vfGByTKtEy0
2NuPSFFCjEGZbTEHakKiUV6tcqQujJt4cJeOLMvTH/lU8M0dyrbSFyTudJaeU1DWy1oVZB2fxSRj
XVkOhLaif2mLMmvijDgj7E2dRyD0Xu4/YfMKNT0XsEtxCncWQxIa9tCA38mFBUsNwwTz1IiMwJ3I
y4qh/80XEUh33k8XETFsaceF+Ig0EGlPMvHjtmVJd1fR8WsIu8AGnL9QwfEINGEvDl/JXLnWPK1V
hncevB0jRtFvK4VHmv/hCfTvTOTev7TlfIW6aVrFSCrMBVChdfpS9hiRD4tX5n3KQj/0MuNN7Mvs
0f6F7SBXPsuvaXKT/OmRx9gFbgISz5OK47C4/WL3kFz6w480/9bswwRf+LzpEI6ZUThRp5TsmpwT
kDvXnxXfnukmJTSzNH+o1KHtFBTZOfG5iddas+mZR5tmI9bK3i+qy7kptSvL6N03LJ4zT8nbbmTb
2+loW9H7RDvODQMtQbzxC/qOa5wdwSk0GTPK8C+N5Bu0cbsEPMTHFtEwB0LrRgo2lyZf1qDd9j2N
GcmaWkqt1VIi0NDntuwLp3rqPzYDU6GUz7YbonlGx/LVpqYOJ/20qAQSvgCh11dR83j9dj+DGvWH
qbxw+JOuMvsMUQfkeBCm/UVAHVwODX0xB6oNqpFTBwT0uXUTyjFdW9/lvvTMbxlvhSm81NcRz73d
qd47BKvoC3BCEzLU+7di31RNSQ80mXFZXox33gl6mLMjAV/V5kIN5Y+Yqz3O4xy0uQp2+hyZr6ZB
gpUXlVRE5FSZxHQhEQ3H1/dFaJmq/fU85VO6KdZgidzV+GNbviyRmahgp8IiTRPB0ncval1AGLe9
XtdnGPuq4KMl6vEpve78rlOSCrUXj9odLvqf3Nwh+go2KV8QK12W9B1ezpubvHXWArh9v8otZcRm
kCAXcVHRyqeQ4+JVcQrh6nCBB4mVepI+3eMh+NMhaVSK35USd70M/9/HBBvu2NbzCYug5Z2IeRGb
FNVB6nQQH9UjcxwYq6Ds7OSPW+MkYCufKB+DtgN3+bYjj8umE9EgEr667lCpSqooBftPb1lXRvay
XIEI3ZfeTwJJCr+bmI3TLdj8rLYLXwbXDftyyQZm2anxzOjczkC2n5tWnWnuCpEacwIGOrkrAeYq
utxGoFRK3vS/P9PJfpGl0O4tNVSCZUv1vEJtR7NGLLhfGwNPjpLD2XzzsAvSa7tIyclH/e29qFdJ
ntJu4DqlWvtKFsCgm0aCe503AipEQOd4IUWsC0OGX3BjuxdKJEFY6hfnoKDZK1DUhUvTEThSZW1S
lyIMhdmvi12Gi6oXulFxG0Cf1BIlWtTHMIOO9rCr6nCwc2iX4FjP+yJbRbIzzITwy/3KtxkjPoDs
0eoWEvrkj3oxz0TyqPwI/qxBPgs3W2bPu8lqFLvnpb4YROyO4XPhZHbd8/GWg9U2RwnLgcSKrKlw
fqvZLYF8xcjESRIXwEOzxeW08PfbtGzW46AT8wPjLQDBgm+pbCG1G9yUhRICA8wYJNQB9yPK/cgp
3dCvcHZALhCapRxRT4f/nHJ2PmDTjEjw612rXfTCeRH4rKqa2WD6bFTtI/b4Jo+hlNSISmXoVCqr
5BKmDdhckq9JjtIyYlIQMfGAjnTOiuB7HCX7DoTfKoX1+jQLpg5YJMLvk52QUU1LLRWhxAPIUGzf
rH2HL9SYkYybtrdXfptBsM91U3MrzYX3G4FrMD5sb2uCDCO5wW+0oYRosRiwt0uhRHhgYBgu03C7
vPLpcT26gjMg/g9xc95KCnGoBFfHCeiVYokvtr0Qxyqt6WMdSc4KB+1cGn7uzrX+fcrxTXtyQuST
GAMgL7FDAZBdEU7NmgsAgdcdkIyKA2xzXrDt051TlEq3LLH1oShdUZHcaUjFMPfUCknPYWOBSyUQ
N7BwUHLbHO1spwDdgdtWYJSG8rzYSot08aQjnsU8sxvUawkMdGdFa7Lt+NUvC95Da2E18CEwXtUP
B89otejaeymBuxBurFP7kZqZzr8IMHTuPmOVBJBFnZwKO4qSNt/sD6wPjyfb5U10rrbA7XV0HLJK
8h+SyBT23zRSRF8ZOdXTBnsZjk6Xt4rnLU8xviJ9+HrdkIgfCHU2ibRhIrHbJzs6HOAy9HtmY29J
+Of3C05g4NZjSVK6p+Sm8AX0Zj6BKlmbH+0v9wtUhqtCK+DXkaDiWcAd0Qms2fE4izmG37BDBJw3
eWsfj3ZMmkDNsED2OOV2LSkhBDlxSp1gdk7M1ZpUW9ufm9JbaBBvi9zKw6xKi/OBke9uutA7mGeh
uK70m6peMLNFIv2VMe0apD4tULS8786zr5hCcwkbeaPECAVFqqswJxS4SO5K3SREN+9nRsiD6MwA
nNl0WHXYWKgFeJ8PcTvFGCYfpMSKLnYH7sFOT+zMvWaUw4Xx1jJyfb1WqJRAnmZ5uMrfSzZNdeGt
I8psSL+3zh6BuKlOpTNYWmkEvD50utinasF5w0mDTQXEPjp0lkKKqVFMxx+kn8ugjQbkJOfb+6df
waIvBmMaWYM3Q8fsVpf2aCJ/SPJIzAdBrAGCw4eDxFOlzF76W0yfXDcnMgqQvmA5UPxdhzIV3TJ9
y1e4qFa+QYWEI5gpyZgEdDy+lyydKXLMAVfYrN2vY8tZbfgHwbGQmps5rfvnuzUyCF1eJtyRaj0l
WYTLH9sBNyM+Mflb1um/VObAcvxMrabfpKU+oFUPuHDgmC49iHwDasbl50J6o6BZuLltLECNYuGW
8kzxLvdLReNM6rCtv9Y/Oth/GzkHMHn5A/hi42f5oW9p5nCos5gFOL66P8PqtKkXFzpJA89jaRH1
djKGG1lZ7zyblaVkdCgQuj11TutbQ9ugL8lkQD73mM1EqLHsoiWpG27hK5UYaMqiwO7TCAcWwEyd
YgIvyjv+ITjjRkoyTMlvrfz9eZH79cnOMY/ySZfEt8txhWJ3RBdVnsNTJz1DieBf+j7ivT2CtT8I
xKXTb+STjb2d5eG/XwmuzpQ7qRVOlsHI9TAKU+VxNZZEUeMSKJlvwDZIRCVEsbuhVyAWkSAWAK6t
gxxljRJuxsD5Gh5VV3Z03oekWRJ/e8XMcl+yksk3fjRWYBoTeBzyOtyCewqWHOVHUdkC8h5ZSyDq
L0xz71Gv5OrqXHtZ2S6kxhmKRx2DYo8KGI/lN+mfbuwI0lTl60Xg/8xmH2sabyc4g7g16qA+tQni
O0Ixde4l3G2VGzKvpgiI517B1DX8iluICzjUH4I8iTcaYKgQeIS6TqEQdtdey5gRn+oS5aT7pWBN
VGjPjSBL0rDB33a7q0vc2ilVUdXpIGflY3vHXd/XbUwrt6FL3UxH6dQksSH50O5flgT1LndbaCS5
ABRK1Hwk0o7feeNNi6dTaczkad+7upH15zp1WB7J+kWT8hL2OOqdPxA4mTHWgIYCgkTfPCAlt9Qf
T8oSvEav1mJ3nlAnrHBkkobQ++ayp++Zggbu6pXVUp0KA78CIAQOu9eH14RGCqvr1NBxc0h7UtG4
h3RpshfEkSUOWS2zISC2a1NsJeLKZ6jEv7uFl5jpFs/PGoyhcHl4RiTCmd3ZcijOEdGazjURlm+D
ipVpZBk1fucL/xvniljQ+0scABwDpYtSrVQ55dymxi7rUTtKwBVhp2SEz7l1k4Ujo0mrZ1TJtcvL
ho5lgIaV8ExqU16iTyPGDul3Dwz60oWUR8CRF1Q8V8XAkIYe5niBS3si85ZDxhyVCcJqafOY24zR
xrtFJZzR+MCElz7v0ukQgKUaTrjUOu4zFTH2/urbQrlDhMbJeN3+AHopIy2vdI54S+hrQL9AgN2g
GdnQAROJCJHF7HQjYQa1+NOm88UXLt3aqfyuAh95LZDMZeMRFfvJjpmQvrC3hm2d1HLNdBLckvk9
N7h1r2KD/jVydFhvDerEiF1SPw6RVHcxkaZ4n6VbZmpYQQwiyXYZ4L10VeFJiji6FKZwLxsRIy8/
WbOV7G1gGhjMHeatvPhsvDVfdEi1oJK5exJbDPwsK1RoUUUlDGugmxrkYiecBp5c2r4aUu7NYgxn
snVWflnLQf50yYyiFeBtlByHoVEK9Asn5mXm2fkxo1CxlojcWn05zSx6LCkTnGVSbRy2Bo7M2WQJ
/pgT5Rt/HPA/P1VEiCRIjgQiiFbQm5FClijOLHnG4B60YgZY7jWgZ1HNvtDQQ+V14fmOEmqBHmSh
rdv04ZI7y5Nh5b9qlLczmK9G3vPo4cZV9NB4fH1uUQj5l5NSmga1YFP0eDdm5vV/cDKNYHOrmHKp
GRXCC9R4xMk2lgHT1KNnXdv0tWNpkQOtHQDgsZvWnHsRnxuYYNP2xSiAwlF8Ohtg799etrohKQZi
AXNhcFXx2Rv68q0h1aJSCGglnSVcsurfBEBvwKu0uWt+HP+wEVNQiCXmDkX9qLvvpfgUuvkEDI/h
PneUcokitIBZurisrZSf29/Z003Gi2UTtubmyeyTWNTr8VeTaFw5dkIEgZ2RX/CJOVuymP71sPKZ
8K7gDy334e54Qad1T/K21OJVESsOw6H4kltu2veGxGB96KJ9NQNakl9tdXDRDJvLCtrTDoi3sp/r
aTVdDZdQJELgtQ/g2lPzj5WWSwzfOOaWYb70fA/EB+BoRvfn8E/inik8rUzn8A8zPFicbXKvzUTx
uWwdHHM+ELaqz5kQSQDJRW+nWLbs1KxEcYZFVSOzAzS3pPfdE8Y/UjuNfV/vFDHkvfT40+TL5c+k
XdeIu7cy6D9EbgJ6ql6A/ejr9mB2P/1Orw8UuaXvfFgnr/gEnZ3SG0s3Rvs9l5sx2IJ+xV4eg7Cf
rUebI0G3l28iv+29x09y9L7ZRbu5I1LEXq7Ly9WQFCP7us/VFWXie3IZR4AWn5s8LuDdO5UhvHKE
x13MN9dMYO7Rv/Ul2opU2TJxE5Lkay/5wTB215w2z5Wbr390sKJc4G0BhTr81mxrPP+ZB+Zhk+nM
V2HWDDg+RdWvAS/VUmdRGjVEVUp9rd+xIdPgIYhCW5FdScqwhFvB26WPq9uqB+dGDCGab+unwY0I
U4iEY+h25ERBIkj0uY6bhITmj2UuYPFJYa2fYk5U45H9Cz/rbFf1v+DWqi97McoRoboSUBzzquGS
DNGYZKk8mEXu6tB9Xi7WmQOQHJAnnz6z7Q5xS/lIIKnJUX0ujXvcw47hYFS8avNoGnXr1InSUIao
840Sx9X9nstnoeX26W0bhalMdJW4bRIYEOOgXQfX8LaYf3KA15Hmqk4X0m3Gq321ztq4dVhkt3H/
zusxjCNYu88jVFbGfX38qqw+iK81+bJwVsVv+aN0C2sVrf7gG/X5Ccc8cTGChwp41NQ057DoSzaO
V29qObOtU0GOXmaveFLPXb6Tx3/WeCRPNgusW7fQ8pe5i0eUOUKo+PN/u6GkZcrNDH8yKhJ5Zv5f
aybFe/9ohEqOUSIgNlcoTp4MthHXmO0rnATPwKPRB+qUWx6A/C+60iWdeb7/YDlnxgyRkSpKWCZU
aBsHI9m+dkJOAabKfqFupJXVMQLWocaF2Wx+NSm5JR+u+vtftpfcBr5I2Kx1TJ/HRX6x+szsrhzW
W66LFcpnjivQVmFVp1t3ZKxjPWReeWaczLf63vDfleb0W9caLrBZFBoR6nUD1Au5OERVzHU=

`pragma protect end_protected
endmodule