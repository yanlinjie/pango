//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//the debug_core module, which is one kind userapp 
//submodule list
//trig_unit
//trigger_condition
//trigger_out
//storage_condition
//storage_qualification
//data_capture_memory
//
module ips_dbc_debug_core_v1_3
 #(
  parameter FLA_VERSION       = 32'h9001F003,
  parameter AREA_SPEED        = 0,	//@IPC int 0,3
  parameter TRIG_PORT_NUM     = 1,	//@IPC int 1,16
  parameter MAX_SEQ_LEVEL     = 1,	//@IPC int 1,16
  parameter EN_TRIG_OUT       = 0,	//@IPC bool
  parameter EN_WINDOWS        = 0,	//@IPC bool
  parameter CLK_EDGE          = 1,	//@IPC enum 0,1
  parameter MEM_STYLE         = 0,	//@IPC enum 0,1,2,3
  parameter DATA_DEPTH        = 9,	//@IPC enum 6,7,8,9,10,11,12,13,14,15,16,17
  parameter EN_STOR_QUAL      = 0,	//@IPC bool
  parameter DATA_SAME_AS_TRIG = 1,	//@IPC bool
  parameter DATA_WIDTH        = 1,	//@IPC int 1,4096
  parameter TRIG0_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG0_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG0_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG0_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG0_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG1_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG1_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG1_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG1_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG1_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG2_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG2_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG2_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG2_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG2_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG3_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG3_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG3_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG3_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG3_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG4_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG4_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG4_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG4_MATCH_TYPE  = 0,	//@IPC  enum 0,1,2,3,4,5
  parameter TRIG4_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG5_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG5_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG5_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG5_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG5_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG6_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG6_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG6_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG6_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG6_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG7_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG7_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG7_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG7_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG7_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG8_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG8_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG8_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG8_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG8_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG9_PORT_WIDTH  = 8,	//@IPC int 1,256
  parameter TRIG9_MATCH_UNIT  = 1,	//@IPC int 1,16
  parameter TRIG9_CNT_WIDTH   = 0,	//@IPC int 0,32
  parameter TRIG9_MATCH_TYPE  = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG9_EXCLUDE     = 0,	//@IPC bool
  parameter TRIG10_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG10_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG10_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG10_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG10_EXCLUDE    = 0,	//@IPC bool
  parameter TRIG11_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG11_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG11_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG11_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG11_EXCLUDE    = 0,	//@IPC bool
  parameter TRIG12_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG12_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG12_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG12_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG12_EXCLUDE    = 0,	//@IPC bool
  parameter TRIG13_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG13_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG13_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG13_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG13_EXCLUDE    = 0,	//@IPC bool
  parameter TRIG14_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG14_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG14_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG14_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG14_EXCLUDE    = 0,	//@IPC bool
  parameter TRIG15_PORT_WIDTH = 8,	//@IPC int 1,256
  parameter TRIG15_MATCH_UNIT = 1,	//@IPC int 1,16
  parameter TRIG15_CNT_WIDTH  = 0,	//@IPC int 0,32
  parameter TRIG15_MATCH_TYPE = 0,	//@IPC enum 0,1,2,3,4,5
  parameter TRIG15_EXCLUDE    = 0,	//@IPC bool

  //   Initial Configuration
  parameter INIT_ENABLE       = 0,  //@IPC int 0,1
  parameter INIT_TRIG_COND    = 0,  //@IPC string @H trigger condition
  parameter INIT_TRIG_OUT     = "3'b000",  //@IPC enum 3'b000,3'b001,3'b010,3'b011,3'b100
  parameter INIT_STOR_TYPE    = 0,  //@IPC string @H
  parameter INIT_STOR_QUAL    = 0,  //@IPC string @H
  parameter INIT_M0_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M1_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M2_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M3_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M4_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M5_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M6_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M7_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M8_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M9_CONFIG    = 0,  //@IPC string @H
  parameter INIT_M10_CONFIG   = 0,  //@IPC string @H
  parameter INIT_M11_CONFIG   = 0,  //@IPC string @H
  parameter INIT_M12_CONFIG   = 0,  //@IPC string @H
  parameter INIT_M13_CONFIG   = 0,  //@IPC string @H
  parameter INIT_M14_CONFIG   = 0,  //@IPC string @H
  parameter INIT_M15_CONFIG   = 0   //@IPC string @H
  
  )(
  //interface with jtag_hub
   input                         drck_in,                  //jtag clock from jtag_hub module.
   input                         hub_tdi,                  //tdi from jtag_hub module.
   input                   [4:0] id_i,                     //identify number from jtag_hub module,indicate select which sub module.    
   input                         capt_i,
   input                         shift_i,
   input                         conf_sel,                 //indicate this debug_core is selected, from jtag_hub module.
   output                        hub_tdo,                  //tdo to jtag_hub module.
  //interface with user logic                          
   input                         clk,                      //the clock from user logic for trigger.
   input                         resetn_i,                 //the hw reset from user logic, it would be used for powerup trig.
   input  [DATA_WIDTH-1:0]       data_i,                   //the sample data from user logic.
   input  [TRIG0_PORT_WIDTH-1:0] trig0_i,                  //the trigger data for path 0, from user logic.
   input  [TRIG1_PORT_WIDTH-1:0] trig1_i,                  //the trigger data for path 1, from user logic.
   input  [TRIG2_PORT_WIDTH-1:0] trig2_i,                  //the trigger data for path 2, from user logic.
   input  [TRIG3_PORT_WIDTH-1:0] trig3_i,                  //the trigger data for path 3, from user logic.
   input  [TRIG4_PORT_WIDTH-1:0] trig4_i,                  //the trigger data for path 4, from user logic.
   input  [TRIG5_PORT_WIDTH-1:0] trig5_i,                  //the trigger data for path 5, from user logic.
   input  [TRIG6_PORT_WIDTH-1:0] trig6_i,                  //the trigger data for path 6, from user logic.   
   input  [TRIG7_PORT_WIDTH-1:0] trig7_i,                  //the trigger data for path 7, from user logic.   
   input  [TRIG8_PORT_WIDTH-1:0] trig8_i,                  //the trigger data for path 8, from user logic.   
   input  [TRIG9_PORT_WIDTH-1:0] trig9_i,                  //the trigger data for path 9, from user logic.
   input [TRIG10_PORT_WIDTH-1:0] trig10_i,                 //the trigger data for path 10, from user logic.
   input [TRIG11_PORT_WIDTH-1:0] trig11_i,                 //the trigger data for path 11, from user logic.
   input [TRIG12_PORT_WIDTH-1:0] trig12_i,                 //the trigger data for path 12, from user logic.
   input [TRIG13_PORT_WIDTH-1:0] trig13_i,                 //the trigger data for path 13, from user logic.
   input [TRIG14_PORT_WIDTH-1:0] trig14_i,                 //the trigger data for path 14, from user logic.   
   input [TRIG15_PORT_WIDTH-1:0] trig15_i,                 //the trigger data for path 15, from user logic.   
   output                        trig_out                  //trigger out signal, to user logic. 
  );
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity", key_keyname="SYNP15_1", key_method="rsa"
`pragma protect key_block
Bu4BPX03qm1+4VYBpGr/I8MmQhBNuRzTZckx41OqIL6s8V6FK15S2qf7pZCtkLAp7adTJiMCF785
xsEd+AdxAK+yb8rmGqs/35hn2S+ZfcrlFb8QcwNh7GDOq1roN8/AueNPSaeqEMsBMZLzme3jF/e9
MQN0ZIb1NfGpPrSIhT2rSYG0shb535mNOJA1J0gyFn4mQbX5bdgenbtWe0+OL/kQxG+AkmTvQSo8
3cZMGe6DTa1g+5gTQzQFd6Wk33nWS+O2Dn2IzhX2awcO86S2HmMjdKiAfbUSfnZkOrAj2UKzCY+N
eVkbo4wrQqD3Uwtfze1j5QMtihq7+BZhHcXVCw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Pango Microsystems", key_keyname="PANGO_V1.1", key_method="rsa"
`pragma protect key_block
mbm9mHGRI1E8tHSEPyYr9ceBOLrLXtc+sJJ9ZhHxkXY8PqY7WaDZrod6DEvny/x5iUw2ocYhITOe
suI31aQau08wt3bl6whew78x1uN/02KFUth7KmdJeQ/OuptLh0D4Sq4BLSuQYWL1HS6YWnesnkY9
k0pRmqJLSguxbJDOTdFpnUwc67Uk3LHO+1ugPo9v+w4NqO85wbA/hFrS/Z8kxMxkHyMu9n3RdCnB
ezQj1MrcsOeK1hzUI1tiEgH0smGunNKmz2i7XtGCOyfiRaA8Y1xSu4iBztmcfUApx+Y1KVjDwJqe
Ji6Q3kdULwp6SPvta/T/utc4xe4v183tU0ivXQ==

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=148288)
`pragma protect data_block
XgxVXawgyBQFtIUgssZxZj1Wtmw1MVYqiCBLIOXdTNo99KPO7rqnVYS8YY6ETx8PZm8LnD2DK6FF
zOFPzC50V6VHHPJVUANBl2TmIG0ESTQR1v8wGrD0MUjbW9hwK53R6zUGFYOVxkYwB/dqaUifpILE
DLZP1yZcpu/6qRuAHSEsaLJ7BShu9AKLH1wnPX9wCa3Z3IH6aU2BbHi/ZEtvHR4FJIzkE46S14lX
zSjAsSxoOHeym0W6k5mhmCQwW2Ht52a0OvMld9S5YcMujnfniRxodpArrZm2RgIhE8PeUY5IS/Py
KldqnpI4+WsPg1RYsjPFdtB+OqDyLtH01Mat3OFlVP6/5mFe4AlPKILYALSPZxf51cfch2teTDQO
Tlgl4puQFo9JNGNoSZcTzad8WuNsfvtW74MOQd++MEmw21bCx0n/B7dygNDdvcj4rHibdrOxr8aR
TcbAzlamkDTQx/ilAbYZHGGQSkBh4RBA4XT2GooNdQBc6RlVP0CA2vQ/ipQgWPMPnRD0gVLG2KfM
18XymJqrIQo/p7Q0owJpQmGT2OAKA8kNOkZHjlnA7U4jbC0pmUta0RT2IKaPovcMeKvuujM+0mLu
zg3aMkh1XbtlXZSQUhsLdtmgiePNYoNLjqfMJ97LbndJTEx3bGeu+sLeBljyDPy+GLHqkrZjXa7T
Wn1aqjRzVr+9aRYdehyAAEoWmf15zxQno5BGXaZScggTrm0e32WkZGXFJfL3r8p/NIlii31H1/cw
zpE3nKo5ntiv4fkjcludLxn8+7Y7hvkGp0XwVce/uAHJ77/YR599UJJ23VY5bOg5wKuLnPrEwS2k
tahDE6x/KOfDlpRntlCQP3azohPTg4i3YGBQY1cEt6YK2AoLTs9AXY4+7hhSa5lbsVPAZucjV1lm
vqCIpmWi6MM0rgR7l+wBBWRdVs3U/F/+CWwuGso3eTtFAv5WBwzlZl9L58M1ePAYdwPy0wICMnZG
3TtfWmzi1s3gH3rheZp+iUnjMo872p6mMwu1nXbmuA26RFyKomAbfK+Dxey/5kmR63+bhS1zJiKJ
PWgE4bGk4Mav8wnzkoTWDs4SFTmDs5b9k1g2UD6/kkVxBbq++qbSLicokHrfe7hJsgPIGHetILmz
JDftGwb0i5cdzzufqaeJS087q8x/3yowFyFKdhk8QiuuFpbeZ1s11TftaRz07+unpmUlW/ScqhrL
V80oUzTXORYw1QNysVWhOhhfbZWEIhznR/Kx8r0p9wWVW2uwruEzd39FjcGwLdsgAKh2R/lU4xUk
9tXu1pLoQvYDzil0aOXsv+dPF1fg2+PFDnGq48rXnAsecfFeQi8DyxLzcGd8mtbwO05Z2rzKbPUA
MkLFUakVuGUuvaZbH+Ottu8WYCAQ/73jZ99r5U06DOGQR06iNldtsy27G3eQzoS31ugCz0FkvVaO
tBLftRT4t6WNP1ITH131enUSWVINoHiWPM2IOrTeHCvf9lid+MQ+FQoh77pjWnQPS8pch7f5SoC/
79wsaspB4gdJnLtQyFtMieV24NbhYdCRfvH1WRTptK3qDchnVSLR2+5wzDk/Zkoi9iDoTLo2Qjal
qwa1J/47LG8KaxDVDl+/bwJj6+F4yIpKhvq01bT57Fgjq3btH/Fz+x+jYx46aKoT0Fs8SssWNV/9
QfCULSETXvPwtYdQrMPCULASrRVg+mvUtedSD9qDVrU8cuvxEpcFARcrkAmho9kqSjQLF8l18Mq7
x1V4/FPJ8+kstRcD4bpxVELoGhRKQT4JA5L/HzlTMHr/OHc+9dKIEA0an+Y485lD4HmOdSAXEHTi
+3VAmBIMrADbuhCJssQVaLHBYem2r5KGX9sjWZASZd2RUapOXVJLpHH2f9RmHfnyeJpCFNpboq8C
WvMIWsa+k/QNn6WiDnN3+4Iv1brT41LK9p7sEH9ifrpe9na2QcdqY/ZQncYbberbd1h0PNEKQgb3
HemMyQqkkuUF7W4AW8ZqqpSOlgbVHx/X9GFHqzH3B5qmxnZJkJlyqOWYQjHW1HGfv2fK8/929edo
ZW5S5W6xXBO5ChHY1nURrjZ5xAqOj/DngSW86Lnw//kdYybqUOZzQNDvXBxFFYjYFo+IXKjAEDuG
L0RLDNxoJwrYLEkmtaMJuAHsQ6kZswQb+sl4UTozdKiHd6Lwyr37NxqMIvz83l8HgbQRQsK/ozKL
4Lc3kzuDk86bBg62W9F23yGZaEQ5StV+2bowoVvcxJ5SP0cAVwrQ07KcPqyF3ekzCOssa4NCIUlv
Kk51z2M3ROu6VsPdR8cPUJY9UrEeUtrR6kJS0qvqPutU6nXk6phzpEOKxFPdplo14e9Om0l/qHQw
mC5RylDM2K4FLP9GS3usyFK2vvN5RQsTDg524GY5MYzOYYP7p6MvcL2MSyLRpeRN6gkhNYa9s9Oj
/kDFnHUiQskT6WTQRQG2GDcXonFYStSSIlw9FTEMzi3CtAUMFBRYv0kFFOMP3G7fPDkZRWMiKzwD
mXNSGcdOop+AGRwT2JQHTeyBYqG6wGYFEFEmSPtGuNnUQvy2TJTnfEIPwuo913g5ff7TdVu3jhIa
OYpibPd49rfkt4kGrMxeEtgXsTjpgSHT2iQCrWXV/G71ef54Idp5ikEoXZaZDLqIvTajtFX2EdvR
T3FYXICF7ELxJgcpURzxA0plCGZJoofyxMD8AOZk9Q53A8jlz8xl7AgyAHRt0htXqwDjSFCLSiDj
jOOKlPTRxzcJq2J9Ol+sbdCg9piVpK6m+bXWen7RmyckfhcqUoaNuC77sYffhdRWcul0iF2fqOXz
mikJPIijWxEv6AlJ5QgNOM4mbjxTmLknfwJ5DxMCVad7bcS1CR8azXZ2GPuP8n/5rCtXhpF0d0uJ
pKhFgpmNU+6/b8uQmHRkScr2K7b39PripZYvjzUc8AKnTHY40Dvihb3ghCJwXvFwsjPuDpFrjxaq
evyd6kb+DQEGO7j7lUU1PcqEZ+zDnuMQkUEJ+pny2zzJjR5F5IqIhU6wiOtlEL6xLGyqwkjOZBv5
Nom0WIxMz2oSDfrt1aJY87GnJrYOcedFg5/2cQQQ38lzk9NhLRARbXNPda7hqh8x+U2cO+CcLnpq
/z41yrZjjBR6EvqDk5NrstNeX6z/Abn6fvYW7fqHGfqR61e4nAOVgZcf/yqlJIQfHWvbfIwNnTW4
iFeFMZohAtcj5vuB1lsM8YlcddCPI48pODgleGBvJr3Om0Z7GvvbKH5BV3upzqveVIF6XDL/kNlW
5oBirt1l7XaEs3JSmgGKBzqMxWF87BROWD2ru0LfJ2Cz0Ij+S1OKTabQgHGBCqYds1QC3Wf1Qz/I
SeZAY6U2bVO1gmcFOHkqrW8uOZ3TLGDCRTmqGkpCR6e54DInsq4CIjO7MMeiB7Utk4r2F0vwJfFx
xqZqBOYLmIlvmhvYqZi6tqwQMMY7hyvNFOodWTrZAcvl5D7u5H2Gj2LXG7L1e5JrjWM7SbbKeRaQ
PGGXNLq0laJZDFTeOoAq3lhmo4hgi/9aPD3RjWdvalU5ri9qyUQW188PTZ7MGAe8Rm1BkExiyUHM
Tor4oY8KWBlOxm1+DgvtpOXX5fTnT5DnXx9OqG6bC1JBBPiIjo17Ej5retrNu9+4hKucTYqbrSqe
lLcatnsJAGTCS/vTliZWKw+KPxqALJcodDyc0Kf48Ld4seyIRd/5hSNbDxItm1ero3Dqs13lDhBz
bIsw68MmfiILT73M2+2ZGQjz6wLFUF1oe3Jha3sOKKTpuRaJKdONJXxTBf4ZAUunR1So3EhYk91n
kgDGY4H9NhKKX2Smrz2dymUMFhKW+1ScujC1/auSLre552YZP9KCUdvqXrflGnir7zYw1eUKNn/H
jux/43rEi+wDCVp9lL75XWJHTj7jb2uAkGBfW2ALUhJXgkA+DN7OThW9BEn5vOMJiKS1InbZ2WC0
HvD6QPknA/Vfjic8TPViA6nV2WPXtSsKF0khOaTyEIUh+M9Ir4CWEMH3g3JY5wALl0+TOerLWuCK
zMmwT9snOp3Z55wTYvm4trL0s8AEKSeAnywd/NrS8dhSpfWJWrR3FEgDcyyK1CmbAu6zvvLmXvAm
GVttrwyRWJsiYo9jThQC622qlHsk6ik8HSXEppvtUiQGFeg4BUqXtl0aAGuTaBU7bELlf/YsH7+O
A7Z6xTNAKMD8zbaZ+RGiOHbM5WlUYyMGH5ivfRHD3Pz4R9pxMK/PcEhZVaZLWX8g/Mx4JBmcrNuK
WNQ/eGgquBurdtEtE7uIEA6wgziXVJQWQ3tTsG8B3yWeYl9wiYMVRD0fVgk17DlddpATDZb+fs+F
BiElXovi90Bot89tNGJp0lKXlhfKFHiuHGYJfDfLN6IgDheNfkEt1MKWv6MhY7YCufWSO0cGDZvz
2AhMRxbAO2+grPS9f7xdGJZhmxT/Fqj9fNg/3WLDNpkV4/A1g4deON3/euV8DyhxB0k/nYE24OCz
n9UWLitZFzznSBfZdzEcX9HTV28zcR+NbpJxLWhUqtFn6oNCSQDrUk9Umwl1HkV27f/nd5arqiNp
MyIYdnJYQwQCgumdl4OpO57oKHII/ZV5SwVvblyf0cjFPLqldPdCt0YmgpoqkReswAoMLhIB36Es
37jnOQOrQKzGeb5b9/TwCMgvbuF31qo/f1lvRtMqhWJVV43HuEaEQR/b5Ka3nPT6k/nAtkBi04SQ
zP6Y96peWguDz1TXPn1/8rPdbk42GmsLGBeI8zIA1A1TCLV8I2iQ+BFnFhiHkNfUswNomiZYl7FR
YZt0IsrFVy0HlppmedkheTnsjKPt2v+/UEjiNYECnXqp9jjik8XOH7sshxatko2zw7r8dnYT/0DL
kMD5Np4Anmx/8RAKkxWQ85NtSdeD4+xFuwIOX2Sq87IQSBpW0+t/R1DZnzPvi5E58yMZw5gARRtD
lVgvswp7c3TCbYAk/ksevHlxcJPvwUVBbZcxIGU+zkhNSTy5Eu04Po4eW9T+rZjgaKvvVjq6Fb7Y
d9g/0KvLzsxSxW/KNi4W7djOcclSfffPBJFRcib7GesRgS8ob8WejicT4+zxGkBsShpnVXcYDNTx
wJc0T8OzQ7gR5lLG5D3HDAlL0R8+J/b2nx9nXgXZaWnHcSxvnEEGjZNIQ28KBD2nV3DEbkRsADWZ
upw3LJTefTClTC/20Jp3jWvy219yC59oz66SeuadArlKEOEkKwM+MUZJOVanOiMv9QZ+p3x2OS1B
yVkosNDur1kNNBGI6+CY7UEmn9ZaQ0MfeOZ6Lrl7JC9UJ3VNdSkvMw9nnJH6pHmR6XjQehUC2Zqc
4nYDs3IIipuL5r4LkoxPjpmePKHnohL6JHArDiOx66got369r40Uq90ry/IuSkfMajvcK9aDKRpO
mBgLi0NTSfKcMSoIcrIPPrWFMJ8u7x9UK7dMzDkTQyVG8k7sAQ/UxJGlHxH82TBDQ7U91/fknwVO
uNngXfTmzu8wbcY/iG7qz0AW+c4/Oa7bfWVtsSD6G06a4KpSTNUUADY+kf81g+zfmfeIhYjNULbP
0zFm3dJ7MiZ6WufnZ6Sk1VL9BeVFi4lSCifleRSZMe1lH087teAxb9mgihE8IT/0CY9SZHkZeR1v
m0SlIXLPv0nZiLULCTiuh1hFPBqSvSv5xm56N2GKFDb3Cc/VuFHE4nkPfvBZ9zlh4XKOmhG9r6Sc
spJMeZvbwF9zmEnad8CEf+sTi/Zh9lg3en+9s+TqsIqjoNkEnwbpXyR/KIqhDJaoh804M+PRYrec
GITau0PaDUphXsGmUrIasu54yZUjuV7vy8bCwkbMN0fT+jR3/CQBDcmZJgrBQv1FSgGe/FBXrM/0
1xQYf3ZqTop7h3TWzwyedgBXgAn/1iXqYNGxAuCsy0NZN4KjFheHQMhqWGbcwOskt/u2s+IbNgoA
rGyL9m46VTSVD0tdKvivRrtD3PPgrKdek+Y0Cf+RIXZJl9zcFNduyYDfim/FmVy5kbcPNetV92E9
ZXLchuOJRfR9WEqWUXbBE+Q7hCyipTF0oDnzzeZh03An3BDIjEt6+2Lornz222TQKsZAQ8vNsd1Y
44MaUnlA7oTwmhKRH4W/GF7WkBrQ5OR20oYLGxvXVz7qe2Mlqt0ySqpTrrhZTmF7dFOc2hj1l1Sm
/tEYTU8Fe83PmcCaK3biEp80K9WKmWXdD9Qwy/+SDt1NWASeaoH3vkxFsCGLDmdc31tB1pLqqP5C
1ggrTfFfKdU4jR91O+MPeHBwkVMmtdUT6k6nhXRmpvnSxt3af6ZJxPzyKCBtfxUOPE8zCSp/FMxj
BXQbh5X9QXRFZEjpW+yHYDFIgQnmEt9NjIzvh3v9qzGEK31lKwfxfSpOKLOeRDYhy8YLBwf2JvNt
OlAHC4vGcQzJ/7okzxhevRPrjFGNxI2mN/oSQt2WmcjdgDV3BOlxzlkA1WgadKicRQuMVOa7JcCS
VWxfUHt6MZK/g+uSm2gtp6SdULE7vzvTWYJp34GWtcdXNTfctIbPqKcn9hM6UemCZDM2jxFpYVVS
uDed3gu1iTCz/ngfv3e3spLPPQUYOejEFAQouc0jfrptouVCHKOmdBEFFGAB7pwyKlJ2ZmRwi9vS
1/608pATNwMCYFBX6TeH/ZVsMLEyYriBszr4laAki1LFiBvP4dOhADYLZtnR/VzHg+/+eZ3Gwkb4
58hRwRf1IlmvdC45GPSNJ2LeCZpyn7cCv2/9bAqRIWSEhjMnAdtyQLZKAXhaGasyNtpZnMHH98Ck
4GPv1kElnKLNFkZAX+/0fd64N5Cv+3SPCiekVuk74vo4IlX0GNqpp6ZF/kVzuAqbEOoLyx6x3Pau
8V+5S+bLcVlBk+KFbj5TpJEbhpvu+HKH8YxYPZM2JTy1ppN1uuT2yy9zsDtqiBgqUzOgfJtmXJBh
EOKXb0xGJ7axHbYIhICg5MOYQCJ3XZZq8o1Vc7XhzFhK3OTvGAts6jdekwPEWWQ5MMZK93zB98+c
irRe00xb3+swoBt34eQtzEOpx46rcrqslO1ZjPiPkcTY84TcXRo5Q611bbIfgXEPnS/H4GdW5Gp4
RLTnl55lbc1GalCPKjd5oJjVw7F9//cu9fdELwCYhrC+H+RDWsus5hBgLPw9V0y4vooeyN0Xj2i5
7yMa0cNR22BUSVgS6/Zub8ab4OTtSqjoBw+YcvDR/CIrn1TAdKBAQekRNhJ5+sPJ67kcoNYV3t+g
431qP3AMY2wvafWoKDuGU1TNACX7QOvZnp2ekWuXk4X3BUnzUN7pQdIG3BlWffMpEzHE9Uzthed5
XiwUH3DngS2UUKsADQ1JVLzI/w2p4A8m99vnipkkMoDyBJvg2ACXNcoLsQx8zgl3UsY0R/qUpz3f
ixOy/lI3r6eJWPFkpAvhrENkw844ouPuyl0q06qfMVg1LvVHioTqMxQ5f1Rw/Zk4ebmjA6BCt/lr
owqlWF0RE8CmWUgNflLrhnegBHcNoOS8kgan7rlhxHn4N3BmOidSv7Pj+IwcIxpK7tSM6cx9zCSm
w5Dfd0xRDAZNLz90dl/+FkWc9m37TiflhAIn6Ldx0ikJZAgSKj8VYz0vId2REXcpqqGiTd1ywLcz
BGeex9wyyLNwdlPWh1OaZQuiYE36cRyF9gLoPrg8tI+TMIg6V68vqDMJ/uhZulAyYI5PW2AtEIJ9
PJQl1SJvp2RtiP9otn3wf1bSDmEhdS1NVhiChGYyhLKTR3mhQts8QclJVZP171nw5KyktOGsNgFI
+cHmMfAcE/oIyQJ6ueuDiO/Y9STIp2/RW1AUkvRcxQ1W8MejCou79YKOn5V7g8hqdoDJQeKV4IwJ
Uf8MUYJKytrDlrg24Dz8idZBoIfcPfDOZBOAL3wyZCeCq/W6MMjYcPT9hIa0alSVJW0Sd6nG0/np
mIZAypQBOX0SmKbryjQ5V2cHnRaBqo0Xodg35CkSZdWotGZv5/OoNf6CSpLPOHqOgrCNYInMeG7U
m7GQwIdCrqs1k8ol5PQk6dWDSsqMAeP0mFpku+H9bPJsRXgj0uEQxvuU2M5HijwZaS6HEmxOFuDR
F9BTcIdzH9jbi2bw7qHdeS0mM7k+ZYaHOkGTICTnuXWadNbcI58bGtsE1kEUcov0KivgB25FYiNQ
VXfK+1biM+Yl4zg1c7oUYP+kgEtdSpKjYs8GheE0jleh6N9Tgs34Myb7IbqduYPTWQWv7+qCK+IE
nXV8Wn4VEruL+xdnE8G5B2IuNHnwSUEr5Oy99srdSxaruFH20qOJBFzLMe/xjpBky7qeJvibCCIV
+E9gxabvsZcDx7QXN2vZmP4wBKHkiuWpvb2ESpqwjPDvArSG1XT6V7pw8nx3R/b/V+32TJbkSasD
OVZV+fAaRpPcY4q/WIY5LS3qy6jFEZKAl72HuNkLgKVEjpOfE1fnjcAU7nvFypc+/hTunrSwkwNX
08aGWqycpwz/5M4z/WBCWsivGANUDwZKYAocxsRew33PXVXbChciIGgHRFNBrePC2suxHmgNTnUN
ujY2Q3+qz4dxU/b3G2SMLvkrrEJYCAyp60U1vPTOzDMFwhsq2EhD7LU+l1O82pofC2wwh/9/UUn+
0SarGGmPH0+i3bmN0zf+uANdYbxjqNHTO8qaAPnVJ1amg8HKA4j+VnA6sNN9lH9zA7gBYZOIt1LH
65MOgPQCkOrmu6Oxyvl25zKeOJCz2YTQK21jUbEdVvJsmyHoJXa3bRuxaTGfB7ZdJeYdrEhTQa1K
46cgV/we5zepuv1IDl7Yq5cv1eA45Av5gRvqH/UtkwgafWPptjNVp40oiTJ0MOIbEbqLLAGQKbqj
cNtvJZJBwSL+/y5RQqBxWgay77PQuw/Vlnl9MSYgW+PWURwrAMUg/cHcb7ISYRePZBAQ1GiDrHB7
yz61bAM3BhXedOoTBClrsXqVmaItPy6IXYprPGsjzeVzQg+qW/gn2vT7ULPa6oezY36LCJmuk2Tw
2F4Uoz3jW8IQft4NDvtnXRK+SSU7KBMACWQ8WAii7/s3NU73zkOBEOMQNF5VulkcmLJTg+9UFHxs
M9J0/V3DiQQfuLBl8xJbTl8WrI5KLlQvRd+akVoOof7jGuTJGqX6UAcZSUrRZIkKj4XYOoUXh6/9
GapmS/IfV+pCia8cSg0MSGzkxQfD2Jhn2D6pm0Rw7JWapf7OryRyqVq2whxF6vqiIXakQ8IhsATS
KCzxStaiZP7NfTV1rUe9uVfjCr5joJt39Qepr4d23tqQiPY7F2T2yFUkCV385yE3v8z5soz1JRzy
FhaITG4pdpfXNM6fMBYRRZT+oZkurcG2yppr6X5NMFg+7YOs5VQYtL1qPXI2m61jdbuzlD1aNfkO
bEY0qKvoKob3Vh7n7OFL9JOXgzJBTaK4z7N3+9YNiOgPmf2Gz/2Tu6690YCBJhEsOfno/Zv8LMU5
ssx6nmWkCh5C7qdkh3b4HtTHRH8dRyWxSySdi7dHBQWeeZ11ColbZ/GRDqA3GAgeUWHYNkAoHkA2
aN3hp4MkNQyNGkCorH7xuzgpBP4kbgR79uPF/GdWcD91phc37nZMPbQ3KXI5vMe2JQddfba147e/
JAHALHuTEh8rOFi400mAyMrzfltPPKQOz7bgKn+sPjhGH/rGhTk3pWuDkkmF0F7m8Jv/+7QGURMi
+zuYrspcUo1dgwDvqRcM3TzebvMiw0uloiyijAReHljW5Cd1pUjxUobuixVFSq5b+Boi3brFu62v
BeeDmFQ4ZYSTZ5xHBoIfNXi6zXXl2Xe+6MJqHtldL9vImWUJuLw/b5BPHLe6r4TKRelk82sK38yU
O5cALf3kgKXhzVYk1vQJ7G561ur0zDgJNGKBYKoPZHah6LhDq1HVp0WXcKjA9Pdx0TCh2xrFSVEm
XsvmL/3r2qFehNPrJkTINYnPZa00p/u5NhnIBLccSS9/ZaX+f466l2iMPQHJCMY88A2RsMgG+nkQ
q9N+JvskLBGvqvls5Mtx3Scir1gaOOrCO29zKiBxo1AqQl5CzZE1A66rgmd4B5vPnj99ymnX/EPW
WEYjnG4CP/XMcVUBKvFJHCPMAvhu3Xzb13GD6CxoejzatKG/ZdSze6mv74duzofXqNJwP4/vJZ/E
yxEc/z28qmDH298KDSvWYFLyizsY/GflxggkE+knobcnFULF5OigiIGr/UB3QH3b3V0OrImpBSlL
iPzOZnx+6xV8ylQd8jCMuS0SThoHOD52cCvlhS7jZSS2DBQvkhgWpn7A3fQeY/3FHC7eVQe3PK+8
xybh3t85XdrywQASOCDCH6IfIlxh5izqNU5H2sA6WzuKldEaLZYvYiyZXODQIsflXTwaenx7N9K/
n6Llv+Xw7RAxxnenfXDYEbNmOhPqNoUcAnzImy2SM+ExNBw1/IwDM6Vqi0LGjcyMAQ9haIFfUqOg
ymX4XXqx7gwhgpG3SwiPo8Xnb+JCdGZGZwMUTT0oifgVNcnj+xdJGZWlylffqbLy5nSXJRYqL1IH
Z92eTXpFq0GmEwjVhY7l9sdAHjTrbeL2g/3muC/ImHse9ShAZyYU1mKtlxNKnyA1Bm907YI16AQ2
ws8mgs0SwhSr6M9avJGa7rkLda9HXJQ9cFTWfOV1g5e+Wg/3Z4O8ly0NZHNL9bSgfGiKPLvhLWDm
TvtaDLXD4aLB1JPw7uovIQFxXZ5fDKVqrRc7UXOq82UNigpZ+jujrmq7VjPZ6rwNqRk9gLWbGCrS
gulygROfCwjY3YaPSLu3OCH8XwC1WXc6E6yLqWe6tASooP+fDNKxXYlBeBVvW5bqbRkyZGJQYJfp
XNRUzIZV64ILyJX1l5iuhjpj1L+9vJVsrYHvf7Xr6u/RQ1fxSVoqk/MeF85DNNCfDMwGB7u/ecZX
+NPu5LpMLUI4biZZtbbXsMYIp7Xi3tX0t5Xio9flcXbz5AGIl4dCzEJFrWFsszku8m22Nt3PAR2w
OWgUmzyQSeSVof7P/inTqXyc1olKWeAkvabsYHAJpv23WF9nTEDCwEBOXaTbSlHIC1icOAqry0RC
VGnsDAE/lZcRptsm84D3RTWX78OPqvOFSNZn+uSY/ucNrvAa5LpmXbljAQ6kDI3RwGgVvpnrfr9G
qj0r2T2Zj+tw0QBYdPCBHa6cY9oXV3EiqbuS88gIMj+Lh8TElPzaAvxZ6Ad0oAun7QFc3UiJ8wlO
acTft9hs9DFly3+0kmHWPNh397bM/SqjtlZydeZGbRbV9iuo2PgmTYjesv5/0iUDgoUOuVhi5oRz
nUPtKK38lsTd5/lQiy2pOzX10pNcZQXOADxmdSzxKG6poCGr62MBJxFCnLr45fG3hs+9/FIFscuB
+amQ8tYx7x7XTMtCXilmTu5DIkBUnidamZJBWw4TGYEn9830eF2lH969ZN0YnBcMVomnKmYpWISr
XMIPST7UvBGLD2frzyxFXgq8jtr+IMRkvUNi/gRQD74ojX729q5lTsPA7hmqoJa8AjSFqY99WaID
9voUKhdoBkQVWdcWCWeAkojT5b1cZY5Vi/gN976SP0qFRJ78QrSe1Wzsc7cKq2m8aGDnc+eTDoaa
YImOJm+bZXOMdnuCMzn19bNMmUijfPHUSiKR0mxHgpvVnZrLNuqTukOryHi2UUZ3X/ZnO80X12Eo
qOzwdLFhe6ioYiUOQiJqu5PL+Kc5DHCzWmG6M1j1whnmfjSkObkp0YQkpHepNcOaATTSXbmSqlyv
m1VB1wqY6a4fn/dDsYR1eewQ1WK4NGyJ5Rhdivt5O/MhP/ANhBonj1p54KPfRovF77yfrBvwsyTw
IquYCau4RHv34H7n2AkYilC6xfVfbSgd8YjO8tWxE2ykC3q4xcAHmtAr9eIkBRNC4aU8PjrZqGpP
NYrluNdhEnzXQpxlAp7bwa+769rltbhXrrN3now5d1xeZjo5QjhA2v3n4cD3dja+bRn2/zJ2jzOD
pBVUxDcYMOnz5jS+k6ppzZqcEMIluZl/GeJ7Fov2j+Cm3ZrO52phH147RVT6JZjvHeXwmuM+ejk1
ZxciJOVuunyiuNpKBTVVYBH6aTfn7Jsb3y6NZpqiJdxA0rcJcmu0zi6H3EKw0/UCr/skEzaNEKx2
WQPpCTzkvLaR77cSQxm2lJhjbGeeDYbh44gLhkgYxzXSnzqmwmv33CDUimLTAL8sbJdFXovlUVUj
6CbNt0/NENAo7Lkv2yN1F2QhIxztKyNe/MCSKE3jNgjOiET2y6I6VX1crLaCheeAB43Og1edaFcg
3KV4A0jsWpt4r0QeX/FCPyHubrc8is8gpu0ebLMkyiHO9yKokOl6/cpZiia/E6Ifn3lAPcaHbjuN
PA/jwmBHfHswwG1QXcVdEpKgioZ9isWEB/QML7EHA5zkfGK7Q2j1X+QzYR/NIbty0NJDVgEkZ2nu
bh7AchlCz2KGgOSKDplQ1U4pUmEUx+HhQkx61DrIzoOy+PKEB7sq8XpoUU4L4jXGz9m07onURwu1
/QUreZZ/Mf8qzBeoB+O74xrgJ57IIggsNof6ws5oT2m2GyLX3Cn5gxw67JKpeD6/PTff5nibP110
ZRvgH/TWvgpnqbcDL1tXojqLXVFFiTxPvJr6QuLcJontGTmISR4Hpbw2QNI1j53q88efjg/nZxaK
xhGKe2cjsKKA6tfQ9wZPPjmYiZj5ZcLgZZv6UytG9nIFf//JE8JZCg+Z6thvdEkYHCyZTkU9bo0S
tGZfVQStYgOOKPBfAkUUO1a3+Ix4wGI+sWcbMCpxMa6M/j4oNTXXZgAdRhe2QAscz0Ny8K28ynrR
IHw7J65WMbSVPINH6Tu28EAvPXm7wquxNx3e3BmJ412GMKT3BTUnRXZM+JIFmRMCVZmJjie6SaOz
Y/DFY7LpLLHCHfvGvKTgOr9A1aJOAmbwbPukX+X/D76XtIsIi5L/6O9Tar3D+OZleJlYwpmu82fP
6vAyr6dOQ53pOyPYpf5rjVbZ6Nr1s2T0HnMF7cJJ17FpGxK9pR9QzEnPXspXs9mroHI6I5Q1bOVj
kooEmaHMPglKzu96Y/jynXSgseoZ89dRWXTAIYdjw83BGBDlid610hoXOxD7YMK6cTce2aYhaF+B
7j1y5Fja8vbGDhwS9cMmtgJIB7RP9btW0bh9UEQTIHFb0cnUnE1E8rGhCtnRevIsCfqN8TXMOY/4
wC6QHXptuTCE2/0eKlhoBHtCr+2xZYi1H9bkPbey5mG9PFI5maEwGqI/Y5yE9S9FU6RQp1E2NnrB
H6X8Kj4VT/VuGIgFdqfLqXjYssoTIlnPRExpbQPSW4hgX8YUoUunDNL8Y378aZHyEs0E6zDkzAvA
8u5iDiucW5OFuX18gwbuqQuzrbq5ho8AUhOd3Ll4A5kBhGdwiVKfeX7dViGI2ENtMZI7d/eoweRn
0xv5y3WvaBS5mCXteK1iR8OspIiJ9GvXMYmAUUZyb1zbcJTWUlgkjyIDDIqj8BsSgV0y5Ypf5YNs
vaZcXP8Ty2VSXGxNh6rJBvpyVcVji3/fL/78MFEUqU8de5lE4IhE2DHWFYfDQihch9e/5I3Zm8de
ctR7VguPV+ynucE13g0E09D7avj+xwybC023YM/Nam3U7bIAnmGVFRpRRO1zwXYo9J+GQ09y9G2n
AtYO17Nxh4q3bRBPaQYaPvYCi8AAyQei0QTbkWrRYWecnyHMQm1Pfe6zrhnIa3DXUUY0NPwmoWIo
WpHMXwk583uP/ptHpbqiIfbzHqf8de6SEBM9xUgUftZDfqtiA2g1DwgY0+DrD6xCQApodleyrypc
o/hKyxb4m/xqJH5hMWS7GQhu0TOJCYl9UzomtVcxQqk634HG/5plny8q6Syf14EZPB2wxbfLNHmg
XVuf9Fo9ePOLmxHe+vUyttZCm/BMRMpO4YfT/x11IjeyuXvU/xW2JmL9ipEkw2+LwumitJ39H+1G
zSB4OBvvqVjTqUcSu+aFNNfRsM6sQJ0aJJkUHAhyFrLqohZEK2bDfb0Tr38AOyUudhtLqj8HyiYv
iU+w26YJbhlH5GhRk/Ij21Rlxhvihqc/7Oys0ZJEi5vc//7Ci7ezZ7qTq4WHlWzdnQFzR59EpEvR
4tzH7wSaNtIWPdO7r/hv4YtUSNW9+rMrO959UEHn7aNscmvrtJNrl2N61DcUb1xYiJio56Ejkvyh
ppnnz+MaGHuCSNUaK0twyt6fOtypJn3MQvrLVSvVBDjH0ONKV7+KbsAzxQ4B/+uZ/B02EFVdqt4e
a7POw9ceLWbDlEpRkqW8cYe1l9V2skarfayjh6aMk5N6uAkgYtE1Wn/0nhSPw3KFrwEq276C4XIg
uScEQaIh3V9j1h7PG83CDNPCEfv6E238wPHc/UeXijpo5BDPDe/mVfgF5Bt/H+utSbxoC+lsydlY
8zeL6QUyHR7hz6UpOwAFHuhZ1e5fbT/slK9CEAuEUEaGR/U2l/a+z599WdBzMFIFt/gSe5X3mqgy
RVdaqvHeLLvgDetxexr25ymA0RUipAGY+6lcYQK6QSeipKCIDEjLXqDReuFr4f3+a0gxFSLw+iqh
bUkSE0vaZys3a0ee+PWqbTfPolGw3NTFy/j0H6sX3wXqdQ07ecPHUtzTqx4apUCSaU+qKtPtYMT8
47rf67a0ssEhh2wJ660rX1ByLyr0Nb9jc8jY7OksgtO3H13Cqy0qwjAcZP25utEoUBw2BNemp0iv
hFQEQu+Wx+k2xMrV6TpH+iZqjndt4Z+aEOvpcQ4Ss4BkaqM4ROlFxECMfrkvTOTa12IFDFqkR+b4
8xIuq8FkM7wIqU8DOLGwPZaRYARD3gBZf/TS+9Sb2+pyqdenqK4LQaT1LTtmf+6iaYQvoTmxlhIe
d6rg4/f1LX6N8cKqVIkxNHDjKHHwlMrJEVf3reqH1rgO3VNh/sfAdWB9Fu9tUkfEiEuSg4ei4x4H
iQvIS9uregRCOap0/Nw2yP7TjiEj2s2sxKgzjqy5O9kgkdctdJZZMB3X5g8B9VK9PtwtrvfBcTKn
r9ypswzncr4lT0/Quu+Axt/aCStCsqPLQHYfe6SP6Kn712EkRHMd/drOIJrzPQfl9I4WwQdLjKny
zg0c8Lx+qW26/Pzo4ZFgQqTscOSp5yPV3FU6D+kgUhu7XUPoBhNYv9lkkunBWedIJLPMaDYdnXVJ
xCz5z7UoCkzLDFbuF6bcrkY+N7VBJ42+ZOV1o/0VGrAf2WIYzrvpOGxucm4SDS9PykKZozofc2Kz
VJLaQTEbhmvT+WaXa3e99dNkDhZs25AnAOaUKxxkL4z6JeaX9WeJN0lclbJVYd6bbx3JiDbKDrss
dHr89KgRmlZjtrSbI0pG+1pKmpiFnC9gLXoddZsAu7H1RIjuJI5w5cH1sSDM44nUbqJxvEX4FA/f
F42RfM4U9GGsMUdxm2//xQ5lmgNhCOvu0EvfMCTMsAmSzzEJBdpZAc3RO8dtxZsscD2G0vSHW40N
yFYU31863qQvVOkXxbeknJeXbLCfSu9i0avBdFGvt5oDwJkoZWRgIgx7dp+vQh0avj3tqupYGOUf
T4pzDf7o88HQNBaL3WkaldaHeOdOY0jv2OfHZhbWzn/G9LC6LW8pfAfEGi2josep4STHRre7fA3p
LusbbJjGT+1QaJ5YMsah4ojlXlH44wGjCTEQQkz2YwNKgAYexrgQvwPlCYAT+R7tnLUG2L5xfFaH
PEys31LfVy86RuqEOsytvLlsgwmL/tEn6dQMNKszOTudTrEujZRNvkYEmC9u5hkzjTZl3qurk2Gx
AtwPdkMjRD9AodJ6nZ6UFBks/4AD5hm+bPN7H5yR7eIYiJnmRyZQ4RBytyOSB7F8/OcRSNCiMjpq
P99PhmFe2zDUmUXA0sGCTXs0mKnnGBPjpq4CisD7KxTQH0ATVd9I5FKWM7hs/cgy3Es+b/kduA7J
xw79lkg9vxxhptsqTtzSuNx/BeMfu3eJyqukmkFEoyDCGe9zqkH83+jvP4Qx4gs7dWb6AK3e0va1
LLXQE8L2bSMussAqeVpSw5mU4XUpnlzbGWMvg1VIz12zjooHWVqXo59+py373HHPkszKV9xnBdw1
yNyXZ0NHxZNbiTViLukPY0dP93mWTbfKpeDwtvde3fPi0W5dRCGi4Nf0yvi5rU78WX5+rcvyqzK0
KnNxO8UGid6Yu/EfadiMWqqZ2yyAXyFNvPUrKoKpBX143cCZgmnGxV0dRjMl34UT/GEQgFWDCWhp
mNahSwdoBOvTNTo4X83Kk379d3tUDpCjrRtEXb11Tbxz7k+7iPLx/jFawd8ykDOINVel6LHX4Pmh
6h1LvHoFiqv8LittkdegN7e2NMQF4mOG9FYa9vAL3A4mG+wvQYtLXRrA7MlolvaCBN0NdEnAbOrP
I/Sxcjqm7BNkwC/AxCK/RMehhdQqtomyC9Uhiit86V5LYzddDAcxpxgEPJvgvmtGw2dXMDJT6pvX
Y2dSH2kM66ciUFh1RvUBwKuCk/XNOtlqtazQbTIs4fNwvUYRHATLM1qjM6ndp8irRHz5xnlHPz/t
MhCtipuGlUQPprKme3MdDKVDT3poQdDW/+DmLaMzwKqpvFc1+3bSytnfBAQmTXg6hgT7hqhOoDF+
E94lEB9b6mEjv5Gnz0mwijPpe/xiF56bng44B54MSZF6N8gg5J/PKQA2JfCqR7+JMgxw+qa5QOnV
sUq+IBlMLr5tT6Eq//8zOzJ+OeD07WD4/qJTBYlaHQuCcbIu/i8bkjvkph43B0Dxtj7EmBbnWJSR
f+NGDOyeOF7kMO3HqJ6AUpdb/ysmFROwHTyDyCgLbiW3ae45rrDj2tMig3oE/ytiVfAmcRb6hDFR
i2e5mconaQUfvuG5UWJTGZ2PYK3SocaU9+G61b8BbVPkVrm8wSrblptMwI+nPjovuYQpWjxGw8y0
d9t+comNOehmTNrZ6A6KxeqW3pnEiRX1i+I/2Ykx8rwDdxMqGn3VFXdPkSXWvq66fHBj5iPadxod
mOayvNrB8xjhHxhtayoDkWvsGRr1TuaOLb37p9mXnCu/S+LcWkw4+bXEBXsb8BgVTNQUQLeA8Z3h
hYPWvS/phFuULT5EBkUoD8/sk2gp1IgtWVCvELGdyTQdzHqjPWQvWl/PZjkrGSkgmMIV5nCUJKht
UVbua5yjJsaV5RmwbA/Muew+KDgKvWx4ZwWMTT2+HWVUTqkkROxKn6/a+0g9Fn6wUKj4tn2XdW9t
P3mwKPX/7xz71dO8jpPxHQPoiuLlrbHLZszd3pXc/FFjDOU6rzMPJ328KnWWHs9ongPXtq1tDw2H
awlslIMpyE8rxtIJ2UjrjChPR2Ir0z+WgR0SyLU4os7RVTGjWvAZ4mKQsQMv0ym0ca4wBhiuen7L
Yh5c2ZbNE70iH1R3aSAywNPTDStXLfhB4lfWPfEvRT7f4gjenIjf17mUHaIT6e3Za9qthFt7u5xT
RtZU1h7cHFkD8nNjfHHJfI2gLQTV/a7/ottet/5B9xKHlkw25Ul9nxQtZMtpcuxZVhLPy4frVj8l
ktGkHrP+fsm6rcB2w9gcU6Yze9+ClpDmVrqHKDuDJcCkXCJr67pawDM5t9xLox+hQALLy+unq/fv
jJm/OP5LX7p0p6nSAJBJusCF1tZaWymSIR3jou+DXMOL/XZHhmlHipgHHRitRvAngz6w7I13rFE5
SPkmOrOvdikmCkN3qf9cnKNit9hp1/VskRFLXoVl3aQOkbowNsSrI3rg7i7+sIxj05py4Jbnipzk
TwG4m5YKfMwlXR51htTq6wPz3/P2tRmucJH7KbPIZKxRfouyKpthvGs6eqKQS5Rs1CIlYJ3BVuiV
aYjBdm5+NjoEI8Rb+CSpeX+40PyLgyJB9MnNEd6q55xcgkcLZ/m9aXDv4umh4UuAA8q5xF27kxMS
Ba1/IMFn6bZJTu5qa//P+W02dthi5fSVl192IiOGCzWF/a83JWUSYZAUnnqIaIfs61ur++lMVE0e
36i/SAwHf3DTOhaXqbUJ1TLYeViddJ5X037SGOM5FYQy8HKYaES+QnU3/TUkquCnaCsv552xSjrL
0pcmd066poNdltb4wHQlzuA6Skim0V85ACXfYzXdSve9FRywjDTbAwoRpQRiRPl272b4gnFGf/xR
qpVULfjE3aH67UpyQdUprSokP1Icc3KVYLgkq6vmlJdaUZ9DucNWS26S4dybUAD3UejG8MoC9ooL
/iuAKMsdCkckgllkdQvjOQk1r4RTpZzbdk8FrG27gLn/CjWYqr8JcjeN4AD7ssEJ1jqbwfbi8YSR
aAdM30z1v8nqX+EgXwytzsRqiJ5Vu6e1eCLCO/CfZzx0w1LUWshaik/Q8mLCf2bb/iwCdtP3gRu5
AvUDdD+9IMzlAriuHkEG5h1vlLJ2naoD8I0yJp4gNjR0pmrJn7H7qVWTE0ouuA6laSqHIp5P004f
EApIOi9LyaprRWEGzfu5bQpiQsS9hilvni9Zhuz0GRhb0ouMApt22HrsvqAW6Gakj2Y0nH33djmy
77Tq+DmJasnklfOrDPQ+FG9BWIP+aBoSL6dFrPTv8VlYGc/16Fs1fKZqgkdMO+KLgjK8/TzHel0r
AvIUso54jWxJSxls7rg88neOyfkwECRevLcZdbV/9OUOLkHjqDpXUVhaPhMgkersPZ1orr3tNgKl
n2TPSyqPl/r70/fjw1cdoSfRhnTWR3/K5PvcHVPlxFY8ywXbPXlbF15SqDwRTtpcSl4sRibLBh1Q
DBI31q4a9yVdnzDL+uOzfUw242MPjM8Rj8nQQPVIxn+8fqu8UuBwEXhsDvYEVc380RDsmzUME4Gc
PEGL2j7lUTj78V/Me0NEB8cOPkR6JpICtD9kJHt01MktGpuOPYen3ERgUwA+472a0dtEwFXJD6H+
0xrIp72xfggaJsyOEglPfrfumvLnCLtngJL5NCZAF7lM67FwqFye8sjQqI6H1uITMaeTRLwJ7Juv
DdqWBdRpva/r/GFMzkn2pxK5KmLoU/yMoKUnSp7+u1ZTBtrZma+8TB6F0Dre6tKaQykTtso2+BBh
/LC2vYjox0dv6ynBbTZBa7ca1q1iqHuk27rZcwJgSJ8Cooy4Fi/NR7CqVW7a34AvwX9pTwE3Qxos
5CkXhVK8q1COrKNa+U+q0Vr4ccIRo0XlaIrvE1YoKv52mkUM2nQ0BY719r8AilftnEmf3Pw8qjCD
58hvsUuH3qTMCO3WLMQJiAxyh+91MA8O5mHUHVKebqBXdlEImPXjta9W42bOoohrw3DpN/GnfvEj
dgnr6GW2tVMpGcMQWRQ7sLZsU5CmNpdFGy2uQMkaRXNiyoutyTSY2iz0Oe6AFSt1E8DRTByuVXn6
5X7SzuQopaJlR4BmQosTTN87U4J3Wph+1QKYMN0VEDmYYh9nYH7gENso9eT4aEp7Av3KJCt0qDn6
AssMQyOpdzy8QD5WKgK/+ar7iP+/PyLWb4o0XqHQxKeiMLVvtklk/vq2clQRnA3ss4HtJd0wx3Sx
2ADgruA6PxVmvmDtX0dSGdbkFU1KOOaWfhlXsuk6F3xFEBz096PoFgams0hMDiFNS2DiXjluSE7U
IVYnlqXO1naQVuIAtT/nDcOy4kD1mtzHrd/PH1hrqYEeBihVwPUvODcN+tRVTZar4V1k9DrehMex
teNkUKle8Lpqo042pbDiz9YnPwJ237dJYfc6jaai3p9UB0PgVafX+JbXHtRuFlg66yzMC/YLRt6/
wxUBU+9lMkXIdGxtR2fCPBjAVMKDNBuo/3kjfSQF1nHd6VwBAV8976l2IBlbfoYxu+jXfHVlCg6q
LwdrRQBZ2eME7PSI8tXC0U2dyE5q+U17Bz4h3lcCYyufrPxYw4LSuFt5VUGBDaT3UQbfaD4N2+Sy
pPKXB7bDrbxmXv/uXt31L1Oll4ZGFBiVBlxk7j6bUxwc6yDeUHP0Qlnerc2tbifj42kRFNXsoR6/
jgN9CbrsuGqCvSSJJ0Vsl/t/f4JQJLN29Mv/j0L5Ywc1dFlqWMUVAlrXbVLSDv8MmRLq5Ey9zwwz
ig0+hAHtk2rCaxdR1Eba6K97QfPyypNEMbEs1WEZAW6lkBXSKH2MTSHVhWho59n2CMVb0eUvFI95
zCadnCXb+tI0uVnMRkUyvPz3mdjt1zzI2uocmKQb+yprapdF3IwTkqUVSBKQSDBoUf1lmY15CRH2
mmy3CO4+AkJn8nlNAXf0Kx+LmahcT8ym8LR1DZCEsJ+aTCcZto8ksnryx+KIMaSYjispxHNF/tXa
0UmAN0LxcTbOCNvBoWIYCoH/CJiXTsmu4mhAnN/PyQJ/LkRXvYsuvgphKNVmcZHInfsgXjU50/Ou
XjjwnNNd2dmUkgQOCSc7ZjTQBTVHQGVWqjs9wKZg4R3EdnURhDcAw1WPtIdWk+m6Yw/LpvuoarEX
9wfrvXT37tZu+skNEH9cO3QhkMbWPhQNP7fjEaOGqTKRx1y9dtd74hBggjQV6vmw7q0s3glG8kis
1ZDodT2cjGP3mU8YP0LP0/hoSYyid7KNSDRwhlPE+2v0ysn9rBmOBkqbEguzyGUQJgJAuMWN4L3y
6femc8mywcEef086UVsYWoUNJLENBXRubOhknYML/Dp8F9JO8LBy0F9qmOyc5zejqEU0W75vdwyD
Vz50HLEEgWzYjJOs4WxbIhj2NxWnctapXjkf01vubU4TbDTCz6fhnTi9PH7UyQeHpj7LuGmd3aXp
5N80caIXLRNo/YVPrn0eNAfBLFT7kvh0Nv81/71Fns+FbEQv7/es07Ochz+hs/6XpyFghpEYdNKW
gw6INJyMIx9a2/Bv6nnAc0VhtSmzCnxRwJsjRWkiPdaXVoGGnkS2JckHVBmkwOkTssT67fZtrGZ/
ndB3+leZjsacg0q1ZIjWi3jcXyoLh/fzOxCzRESWyxmSBhoFu9USlw66sSR99pPkrVGFJtvmDQdg
vphHl3+g2nYY9/kB+duqBVJFRIjAcOKMGUa7TCPoxJkajZeVgCszy0Zak6rp75d/0Yt6YX5T+2Le
Br4ckXCVnNjyHeuqfhq1BQZnUOqQfHk9c9vslHEPYRD15ftj/fS3OT7pNS0Y+NPNsKofR3X5CCx4
7B68pVBx3IvVIeXOzhN+Ddvxc9OFF5xQBGVHjnyzDEoQ4MonyFgAu1Rax9pm5yfjX1AQzdXnzjaG
BdphRJY99SV4msjGhzOatURV2xrvbaaZMzu1zWAaBEsD2QKODoce/bNhedgrFClfO7OgsBurgcKg
IWyf6Dj2BbVUKpRiLC+xc9COyXpO/PysD0xy8CV65WJSqNzpI709ryhZrTmrMVKmlFpa45KnubQa
AM/zxLDy2ywXKj3P575L7ax1sjR4Im/YCSf8rdpdDiLxJgp3UkaVVoTzONwWJ2UtmCiptNpRbZSZ
d01ltk4uGYZRb8+A/UOTMCcty0K7x00VZigKUMTRTI+s3U8mV5z1oqRg9ootKcm8SS2l/a4dcHt7
C1eMGHJVb7oliCG2cjLVLCFJIC5cTiFo64LM2iHjbF5ZXB4K6Pcstyf/BPR/p0CFJ8TcHjIV9RYt
PmhUEVM++bU+9Q65mciDkJw0FJTH+7xb6XTikdbes8KwQ3MrkK+Z0rynl9i8YZ/CY7o/rlYbTe3O
L4jea2tn2whABeCzj2JSxKhEoAPZ8TN9MlHc+hF5enb8HLwWU2c3RD6xEfO1U2OJCUo8hz/Q1Kn5
aubQIyjlwVlqoBUDt0D80gtoq9iP5XalyEdD1O6qdzki8kZSirqyCyLCbNtnNpvsIdk7mcmqNl4C
8RQ9I0SDhbxQk1FJRSi5I4nZSeqlXmlydZMMy6rYx7t3ZirAb+aSOEdhN2V0XOoTu6HlxDQKNZNP
Ag25Q2mnmXzrHsJ5X63G7kKIGrPLeglPm7CUrpYpjcjEp2D/xIHIyBMWqc1w781JdU48/v7dKEu3
MiyOK8x01ZHhipYhaV++nVkSyNWp+t8aNylii2FMOAzFtwVONWc1aRBcGWqN3t4g4qvggZd3R4uc
b/85k5O3BhqfEcyUVGY/U9QylGV2tdzxSg3YrUov2KbYkyaCXEqsV4CzDRD66BPuPAqAFDqTiYSE
zCcnAkz45DxACjS5wTfms0F7UUa4bhGcWbKKyT3UL/bn0JZUrmcEmFoJajc5DV51/3/MmqWFwEBc
UTxCGQ1xOn3OHfGD0G25rqGZyyJCWn3OmwRJFO3yiawNV0lL7pxBqSYTgSjlkWLM5DR4vr1OpKUa
oIsBbrW2wGUgvvWS/8vV/2xUmi+zoFFaN+GmY3i2/9CZBdr4zgfuqAHhPkhk1m2+REeN2ZPUawU0
xUzxDiCV4nNenJ1VzYP0P7wLoEUszL7BWYBm3n6AXHOemWgjSDPAKIsBWcZ/wbFjbc09E4Fs7QsN
Pbr88gv0Q+u1gTK6s7bRWovOEexRy/KE8+2DJnso5kU3fFgR1YNRUV3j/CEiBFmkF0ta8f7NdvpI
mtpin4dIqAI3vdcdkxNA/YybqQlL6D6LGqLxzwL8pQFO8XE+IHKHzo65LLeszBvW0ex+CGhEPQNa
nmHnWPEsBwE6Hw00xRgoz4i96bNogJKHb3BF8gPvTlUOYm4lJtUIRuqD3fM5f3o9FKbMLEoIY52u
JphoJRGRQVyxDNuNzMkpuBW34jYf3lCHNqLp86gDgoi98PJRnM7nLZvtRLrOSfC6QVV3JXZ6bNSZ
cfUJ1+/HLM3Gq19JloUyu1vnguSri9dwU2/eRtYFI2DxwahF1/beUkGkJ2XGoZrtLVq/yFg21OfA
NbAUdP6MjcZuiRgSU4OMrQ5KutzGa+YAQvFZ1ERTw0oo96QUpkySuSVG7L9lqbv3fU2HdCWY4qfW
Nqk1rP7hENx0Sm3jTj3v0vDup0OzCxJPzfX7Imp/cLLSqhg2IVwXxMcIf5LWkg+QDgJxQ/TP7NCe
4TEYpjMo1wTMoR3eU3W4qIqi/mac24z24t3EdHEJDatQiwEtoiXn8hu3zTf/pz9b1cIcYm1ADxXS
RUWlDXkjXeeZeSsQ0xASoKVzqHCTwvEK+36VCBqRi+YH8/ARd9iOw5V8ubG0ZE5j51OG7TQO0GjR
3X4Xi0YAD6DYSlx4U3J0Mr6yQe28OkS55eQzmOltivzuptYRCXJrksaLUBP//J3KKsj63CSaEjpr
XaOn+FW725UM/RiaeCTZ6qlPZ3ZWMLFRvwKGm6uMFD6fmeSRmro+oX8kDGAWzrmTDGN3YWgm/TzP
yZFYL1UunEthqMd8sInHOEWaXmEK+tT+A4+N1Dxr5SlX42DdR/eu2zY+Xd0PeVMhqY5lILDEbzcQ
GO0KEqEnm+WGVWfdauMEx/AivKfm5wBvd7ZQPdufuISWy2JTA/RxM/NorGD9YqGb/+N5XhaMMWCb
Gw0H0K15rzLcdlw5FnBdmizRdSTQEmoKIzM2nzlfx8iL/P214TTmjECL997D3M2iBtDEMaG3Xdc7
DlT7XKZ3btYjk3795HhkLwWCk+V4Zqxdzft7hAFVoainQS+sESoVXI/+1Tqcx8P22kppkpIuRQa7
Q1l9qSOS0omu1wKY+p6bYLloxwZBeYmiul2Sqt4q6q1SKt1LxNUxuvclj77rbilvxW8Gomvnh4DS
n826EQkhSPHZXMpUHfcRjWbHjDocHFnmH6uv0di5dGiEib17SIKvi8dwqjGDAelx+8iOvVyncD96
bWsy40ZA7S82j6Xa6DT6VSjNJERRJ690H+Ea1uxWP+0l2wBErnuMUaxYtQ6MgQKfUPQ2Z4OCmoOS
T+Gu1k8DuPiKSKBtP2KBly/s+9yWkl1QaU8tjAy+EDEInZSn40hD9JHMDusRVDluYrlp7CoWD+z7
XtGJbc4VXsgrrnVLe/2UHQ58Fi8I1Aqq0Ybk7RMCLSRhqDZ/mrw32ajllqfk7uqIKFDTRpbcRiNT
UX54bZ/vXp5x2hrnbNt0OCBX5pTPL7mrYoo8OQW5q4x2QmuFilXPlYoW4VL+1oefnNpaN7bkRQuY
nelqTT0X2KhhYLZ/n7pN5K4MhgiIboonD+ZKC+LzNwb7vzGxp9d3oqwIFsusR0iyx9OpsAooWOvC
GbS/zonTE2VH4mh3Qsrxmk1L3DfaFuvrM2G9HG2nGF1/nwc7AF1vpuzJgxukXdFALy5LP+ua2lLz
ermvHCcP5C96EvPvMFeVg5zBQJqOTzciMDhr6mc7AlDh9/T7bz5YsyPdGhnW00UpVK4dbSSv04Jh
KGdmvk1puPZndeBMr3aJFjHpVEA7HLFm9F7sMoNFhp9m0AC8+iK6Ha5Rz5bkAa+vyPNayIFMQEq7
3UIUT4uGIuxhmukomMA4U09NT0q7k5ieBnX4xbfblA5yWooGTwbVCc1HwWtbnNhUjC5eeVmwN+wT
YfuvBvo86xuzxLvXJUYa5P7gXtS7gWAKSvzS+sLO8jUaujlRfMdijZZEEBYRamByoMZMA3Njyj5O
dKNRgP0OdqXy0KP5US+VYPjOUxCi1JG0/jJp13OSkVsdF5rga2RoKuulK1zrPgT6uOHmSX6AUK3r
GQoDCoE9oGNApyReVudvr08A/KUaWu4IU8T282EC3lXatlBZRG2vkQj7PNTqtAwc+cH5LkNq/V0K
RgFLeO8weLnARIuKbjnxxORm7wiaSxbPpmX+uRqvxRl37tcXwkBxJ6b3ZbctLgC5Al+sp3RwWJTq
cSVeatuMT8nJJUtbiDL1yuIDqXMslcnjo6WLZN5Xk1J6x0hX9hpM5Up0Zrkv65ouuA3Dt2g+17rA
3u3X/4xMkj/xVxaPpFTYfkM7j+NnuR9yDUTrM3gqHZeJjgRAq63OYdqyyAuOj6MLFn1I2MizYnPE
+rQ1yIdF7TznJsxJ5P0zl2mQ+pGX9Z7aoZhQ3Ykbnqjuh6ZH1I3OsxLAy/NxDHfj2G+1R6eEajF/
1uYol//NdbKTwju5eweDaeckHfQ8Xqi5v06N1Ohg+MFyLDFx3z4Lqj+raly9kMJUG8XouTKBqGSY
vpw90smeJZQMDTq95cW9xXDCtUHloazJuB9NeLz4TrQ8OtURpRdJJXD9sPn0aCsI0sylwItuQSYa
ykTwWR87n3t4dqN2DDlLLsyVvcby5/9LZHf2DfYDRxtAYpNqItDNPRSNdWZIKsW2k1CXUkSm2O/x
vOqhRhyJyM7/32mKWb0ov7rC6F3CNnZvDIJu0gw2McDVWAUl+/eBoFEzYiB8KzzQY8Z13rcJi+9t
Z9M24AHaHRjkBSifICvhK9iuF1/L0CPoFiLXkZ1o//PrOJAHcdEPjLRpn/TeaLdmc53GFp5qYjf/
IExnkiKYv0pglyyGpaRqpjDIyiTyWljQdl8RTwjpebKBJns++au7emYEwUGy4hbM39YK0EltUHsA
ouNgNakoDzcvX4WI/r7jGAjpIqGn6k5GIDO8OLXC3uRs4epY2DxUFsC/UMy2Ehn/m72Lt/W45LDu
nRfNePrFE9xmOOtoWdaM+hYc1tx01ICw6PykhvmBEU3cGxnTZB/OoE7RsI4hXWe26q8OFkVsIu7R
YONV8MeTBk0kfn6hOCBTQj2pv3BVB0OvSanMHwJrIgM5Yy1G7ICtXvseD61ewen+f5bRaJyl/AIW
wlPruUXaZFNz70NF01p8jY+01/3KhbQ9TuqjUpPNzyd0NQHAlDtgCv3hNrx358N1Yr/JcogNyyTY
cRRJxDfqDIjqcc/RV2WTnQnqNYqehp6Sy28g/g39mdw1iErgkYcMc4aNmNKywzlDwGaDLx92Ck6Z
rYHIIe7nN6djzH4jPOvpssMrgOmQ8JR1Pg0L24Se6FhhEy5yF/TeRMsJeHlOFTniVjvyVUszYi6e
a5kDihAEswFw/vafz3mkQ1El/3kyVCzQC32UTjTZ7MKt4IsNeEZnUixwzWi3rJwMwCMPkBEs/dGc
asuUUakFlCnOdh8X4AsKwZiehHjSOY27ht6QDc5t4YPIE/rAPKvF2oVQZ/WDIGbJjU2DtnFdZrPp
vjMUzJ8nenWbHgR0tHRXbSCbfLbb5mp2Z8BwJg6iJisOEno0QOwgQXOki+eASMbAS397yZC0DUmL
5rKGz4OaQ7H5z2MAgWGLn5V6/j+nzAm5isc2qQC/XJf+lW1wzY1PxrqszVfcG4P+0sYBPGRp+uIi
N6RiS+auzRcZhYfBpis21NcHjovndfI2e2icfWYKC3FWFiqqBTCbiNEEu/yfhDQE9dFPa/1Y4VHU
k8qbCLMgI115NOV4OxWnV0T3A9Q3c7+69TJpzL7pJqrS1hCDWVj0HWitYZEVaEt+ZIv+IJAFJB5u
qFiDWnPLMCjrm0ha9v/Ncir2VFlRm+GkSwRowdTvrGMaodvdi+HBd1ZQKzOkP+kXvXi5qdEHduXl
6kJsplVVbUtlca4g8wlHtCwPfU5bByeYE4ZImHpKssiFLm0oJBIvrXoAzcw4KNcDV9oifM8uM1sc
pAF1AR48nH+KGgy3ih5pt2721x/e7NW0dINDn8y3Qxd2eOKc40h47SLAbnIVtskw5JyYpPGe9uGe
Hh/jlS+sLl3vTl+mnciO8VXxS7IcLnYr6H5TGSk1xEK0LwbjtVHYYU/nrQyAunZOj529ALAYNgOv
c09BJEsVzNwnSbzSP2YFYVEpYCEU84hYD3iRbihTRVMHcDWnLfkkGTHv5tQ6EN2eC+jZwOizuXZg
8xcS7ee6xxaDtNkP4szUgbcQJhyCd2T84Excf6d8CfDC9VIdkvlxwR4PCeUo9SXioWEijEKmrz4S
Nii6dRj8vMmO+AFm6C9LXCS0lunbfawKQkyeOobrHjwPdl+22D5cHxmtqFvbNRI6Uapdd3HfPYyc
wusqECmpIAdDA6K0bDz4N9PNeFfE6YlSo6q4/hzMn7IpJd8zASxXWCq1viXtJ1MeBf2lnpvxskwm
+vdmQ08yC391hmzd51PLr0joNkvvWSWYe3ycU+0lhJYxEx0iThRr1seYtH+BEoizBa3tZfDGAcWF
yGQgaSzn6VirNfJEG7n5pSykTHhF3f3sYZUh97PYp8I7vzeVUILlKtPZZSHgOFbKx5+yD1OYJaNw
cZDjbEV45ONa8T0WPp1yWiBahuPkuooLzsFhuO5WwhRfxgk0jcVYxoZ4xzpNxJ5i4x8LTFfwiGFG
o7Y5WubcSFFR1gLDaeWKTOItUSxhggejpCzLr0UB9cv7y6lrM8M8r273lR9L5Mun1M/TM8UWglwD
Th4ZT/DrpHfGIEp5QJDSoFEmk2+eG/Kcl2xv1PYEWtyGDzrOpIy7viT2ZhlHahssPBJKoNcrcFMN
jPsp1eS5FLWDY4yKXJVqVdXjqBn0xAQgWnZ/0EHTJtzKYwnntebMIrPmKTjPvc9MYLCWIGsPBEFR
kTneM+wdwWuTxXSbMUX0iGHdNQhBR/ydExJM2jUNXfgCkijmAuCFJibo25ZmKaEYIjIk2Jm5ZX7g
5OoTwDx09/fDAlQoy5bxQXlYU0VtGc6vLffqAc6300mgImn8Y/vO2LLOCe0ubVW2GV2B3AWyXe/9
SgkVFXfyG6NZgm+0hRimzky6qXBlZUvj+nBrCWtv7llFIq6+sD6BGWFPCTYUpUwxOdTy78JEYSms
v0fEIaxvJHZrIGiutx4OeAqPDXWg9ozSvYlcfsMqfw+Q9H+ggu75y0CaZ0YLGkiPqgZ6+RbVWO/0
UdA5ej/3BslUkV0raky2mHyDeaXMXuMTrB/8fExW6GHdU/AQtJPm7iUzuGlcOuOGJ5gXx78h8m67
FON/xjNy/yK6hUvsoyK3jfQIfrl+XZSV3EroAyIVn1nDRBhrrTeW+d/Y06snr2zV+sI41eLJ6aV+
acVFCb6iihPw098O7FP6vIaJ3QrGZJiyg8aFxSG8h/Gp5bvj/2QHDddUtdVLL3VFqNWckfGCgTh9
3aVa8EwZ/rf/vNyABqGyErHr1RENlkyy1W+YwHQ8vSrSc8bEGbnYdhkSEDGoGrCeZlkufxFYgpf+
0ZhlSVERylBRzwXNhCiQzsXr0HAG+TFa3uFjE38AWRQEV9XMRN2hdZ8W6W2IUzgfyl3WhSujP13L
e9Ap3gdKLW2/auccY3aToyeqcB8kYluSGAgBxOPRXVR9h3fONxIQxMPOlcMNFIp9MaqhCCq0KhS7
PsNltTLBqA/GzfhO/900Ii+kLAFchl1NlJaMIJ4JKdbB7LaALt+Q7ML8nCOkDfv0fTSF8p1fAD4U
8TpQ++v5LEJnxZYcttkaEOSLsv0Y28ll3Cpianf3zk6d0rvAPdxBeieqs9HEKkmcQV/oCrbSHZEA
kIwUD70zFW0J887seFW9n95UuhVIyROehkakLkNfKc6hbixy1QoD2Tf8D05hAWyg6R1BkGwmj122
ylUo/8JpUvg/s2GFw93hwoEZsW9lL/RHVqnclL45H0EjKnvJvWUnG9kDCVrHtqHLu/ts19Fa6aST
sOgHc/XSC8HO/gMrpfgKhZa4zzJcXrYaDT8iTqHDp9tijTBm9oiayPjmPqxLP9ydgkGI7MG+0oBu
WRVoQEQNExtmpGgt2gf3b0H8WEob8o942o3iEo3iLVPf/oxMCBVkiDIUVQBed7nPC9e9y2B8nuEA
cwd9n6EwCbJm4pAiCnQjzFQCx/3e6SrJdHWmIUsEd6xMO9Cr7QTnt5jMFnqKQ3JYCfCyyLnvm3mj
j5DapX+M7UCuZglAJersxxYMGdKVXr9vYA7hcUxKZXMnGSeJrvAo211ySbnsiffjV7jilYq/9dFG
1NyzUhRf3bf273e9414LfqCDDPQVKepfPiYtwZApwRNQKo12C4nIHS22aJw/euMDONv/O8uqXgzu
YMe4dQ62szk3mTnNc0ZO9JQhKY0J82pKtHwUoBdi8xBYcIjjYqB7yWBE0HRxNkQuM4GdPXXt4iAW
1ZIqpJOxBzaUr+xdGkclkb12jaW6xkyrE2r+NR0WHEVeeWzC0z489ZxwtUeERPHtPqy8B5qx24an
f2/PMWSQbWXxTpJccvuG7yQSWLkoKMqOdkmcEuapmsUmB1zQ7T9vS20QYZuhC7PSd8LADPiDXiBU
6gwwfl4JGTydgSDgq05okzDIilN0dGYTtQhAd9HmxEq1+bhbsrti6xIOvrE2Xdk3SJz6xHrmpuwE
zSA9G40ztF9ytNThqCQmXqn+raB3Vb3hHsl4+Z204lg6c/dpkVDlRSsNQ3j5vrbtFvsmYV57Ftuy
mOC9QmPELwKTF27Nj38/tUanWCGdAst94XF1iZSogvQLG1FgArCxks1CobuEAkDO9z+moIV+xD7T
9FXXSvcTGg4gmtEcLZtW3aJbVR9+d9FS+DafouxNTD4N2TvgO6OL5/mjS8DH+d/v2RMO2xUzbUVF
QWEB8vvhhKUzqfLzehBoaAPJY6i89D9x0LhwmFC3wQVl2a5b0C/6ki3tZptULSBPQjAwF8kU2vW+
0X0SB0pMIdhkzEOBEZRGw270yBncms6Qpg0/izea1Zn1bnplz12rJA7goe7HDZ3zUQgb/Y/jaFRX
KXnJkNZnuxIB/7pg3w3OFPvzC/CHXj3Hfyz/vYwquYP4m5CxSSdHmpOg62mSju8oQP0Ys9OegKgU
Jxa16UPCRywMpcVV+mlADPWUrvgjIhCvavWUTsaz+0WbdhgXltqELzeTcXLCMiPkoa7JK0h5aE+Z
g5ays7UDq0DaUPFJS/uWbCV2XMXt9riYOaULDXCazFEzL6yya84KmY7rJDVK8dvFeLTmQXLdRodo
mqYFiEPKOKtGl0OYT37DQkpg9GhvEJvPCpNAKrBDTAY/w0nfphkJAZ8S3hXa2pEGKQ/d8AZSP49G
XInFMRTVP4Hsm5ejdUilO/CQ/3Je7W3+NkngWhNgtgQy24fKadxID9zxj8dnq+k+kTqyrB06dDZs
NHkU8R+kkSeBQK5TS5AcxYQzmKQ5gm0BxyfTmTELJ4VyuqK9yZ17rf6/+QJw/dFDLx8E5tS+y1ru
b96Hx+gkgFT0bY/az+vZwyPW5TxTkgXlbAPwiPEABfPH2j1fY03Zoz4B8ovn8AafmXDoqabDfktU
svLzJc0v5c9VMTjxQQHCX31Htt2QRZmxJf7cPgWJxUhVplQL2Ig8Jt+sfeMBDo5Zxtsx2DKVK7Q2
72l3Z+lh01HRK5cTH0+CYNzJhwigm7+MlJy1Kyr2/HJRAQE+bImqDwKhq20BMRam0rXqG2J2GWUz
V0G0CL3HD1ENAKbBPDkCeIhbyufsy5eH0GYadfCe6PXo/X5m4Cc24ifu8QAjAjQkIZ7TQOsuOWCj
1HQ98SIRMqaicroGofM7RJ/t/jL+8zAjTzKGahWC8A9sH7cRHxWONPoCiX51PFdLzE28T+7kKbQ7
JuDs/IQhlecMpOJwWMcVOdrn02UR0Ii18PuRAXC75LaZ+5ZYKMUMdZnSmUqgGxHSDbMpsgiH7WpH
W5DfyNG9j4osnOwV32ytDLnAYnvot/fPyFTiqBJ8dsz6MSgbQIG/j1psg4spvxtY0zKBLKi5zckX
bC6/zYHvNPT0feF+/rEuvkuBOOndc3TGnao2rRLMCvua1zPx4ccqm4eEXUZcSmCdJ4Yp13+PJZTw
LOvFRwBXt3OGRqPxZlDg/rP/eZKYuVgDUj+v/RhetgJJ338xeGRQ+L5C8ZlLBdEiL7okz99IyI5N
M/Uq9njt6a8SKEqqXKdodo+Tcu7rrTQpWm3ec7DpY25QMt0AARj5nIumjB5g+8PDyLgqBEw5Tpgg
5+PPJ4jMOIam6N/RzFm8VJ4LTNz+5JYvWTQ1pbOxxHQWNGCsympX8Fze6hO5P5WhIWijCJNyk1rW
erqc0lCNXlT4d863r7gVyORmu4UBf62Kdoyco4mKWQMWc/Qmum9UqAFoZAxMf9t/dPtqZ4XYGcep
G/2qKr66W62SlQb4J+yce+J3cJ5EST1pw+BFrFIAn6m8f1jN81MwEn1bFgJU73XfJc7EKnQECXRr
1TZnZpZjGs5Ul003zPMvJskyB2VaMgWEDr564gQlfeu5bmrfi6CgSBcUEKXGeJPsyE1Z9Q4ymvYn
QgJAiB0f/jmHtj6w16675Gz7FX5IRoyuxZtezRRyQ+0M+dXvYnMcr2Rdw+cGFpthvQ8wDK0DUvdY
9hdmm0/INvYonkJWtOLp9t8g5xE+B/kkbv3l6BW8f5IhjoV4PeM2FlYrJ8rnDFdu+EQ+x6NojeHY
2vDGYdaKlTu4Vm7PEuJKlAIG6cXLC2pBkvgeTIh+XmJt6QtZORFgn6rCz65jOdZo3SG34Tm1jQVZ
X8OsKy1ohmmHKlfpyZIQaDWGA5UK5xwUl9mO6aRRRNAibXH/P5yBb6ZfLb7bI4hHEH1vVmmvXqQO
5YtFMb6c9sBJtrghshc3mFv6C3rhafM0gUDRLm3Lcl4rSYBOm3tpk9RzZVYH2kNsdMbps4yam1Xt
KyK3MQPiMTYxY9Szs25NT3+JnsW152p3w2popw2kRjkLyAdfYhsOXi3S5fZr/xDSOT6v88LkJwGx
y4rrL8QfB5hVCZoM1AtSomf/Qjal6b3bZnYAen7HB74BSY0OOIf/AhxYU+5PJgZXgoy9KfSdv0VM
Rf1JOOtkPZhAHxlyox0RkP5jQbPseqvF6UtsDyzBVARvgRHWGCIbZ3tOLBE5DKQlSCakaXCiP3Fo
Bz6ztHIhdgH0JhabcLCRT5V4ismn5LlBJU+wUkisvJQpUWbN5EyU5MJ772BEaKPynjJ0/K5RZLmh
uAn6zzoZVDcpvMSK1gaYThLP+BWvjxSNDzOMEhfoO5UqX3JHYeknDrTKkWCWBK9sYPgcDAJ43Y1s
HrpvrhGo21I8BnjN5XWSORM5ZcK1PxDQtrbEIXzB2O9HUkHqTFAiJWkVkwhvHm08tTbQnSKG0F72
JtQDpcwBRMCmkTFa4ltUwKVsEoMwlg0htV8d9p/aTdi/tuuUcvyCupphzM4U8TNtlh66K3c+hLGB
UwV3ZsZHYRAlRBfJ6EGXMSUqiiiQW0M2rValxePX+DFext9fVul+DcgGBhSxrkBO0cKD/k7GbLcj
jx+HdIYtyB+Nzf9CU69xxXUwF/8K9P5wOymimK1saCceW8SnZeI7QJue5z4X/LfcwGFOzqJ6u9yD
QmW4oG21je17IA+xVj4ms8d5O+v2rrLOWnuCbubsm1qx9+2x5jR8EuBCEkh0NkNsmrPfwhztl0P+
of3a4sF2ps3w7Vrzic2h9Aw4yJjABKOG56B8hZXCq7IjOkzt1idiAvl1W+EP3NkeTtLMul3htP3c
1Oq/75Sc8wYVL5fEGaNzhTUMggxe27NCKl2m4FLp7ssbYREikVyriabVjHMuGEAc+TgU6sWRuwzR
W0Oth9x50qbgN3HWSZTsIhjwKnPRsT78yEFhmJdNd8t6q9mMEozBnP79DB6vKl1TlJOB57LKb96H
/Gu9HSsx0csyc1srjkp80W2ghzh5RDpvqSMKYdj0b8r28S9wxpch5D6XKpDnRCKsuBt7NZOc+7nG
JBQvkCCcpAhY3e0yLSfT9Ha9cNRWCA0FMbFfaWiU1VwDjX+pR6oJ8Bfd8OmUEQmYf/REgNNiA6TV
a1sHVFWj26Tu0WOwnPj6wfKVQE1VB7PZKVjwfDF//IpICG+9ojq5yOltc7CmSHxFNIw4sf8q9DxJ
J7pNUOGZGGAXFniJSWr3vpLYvc3VivF4C7oWgRsyGqFO9gAuQyxpbSV0vGvvVzwCO/YqrnlkCn8b
9RJ3B9cyW94QEpSets0LKK5u3ioMK82SlYFbJM/WKFBMTLALSNeNhgndgS9yVI2TiE0fD/3eIYFm
FIMU3jUr9H9W1Gsu1k+s49pcycZRoPzskwsCzezc+L9MGPXD9RL63DprN4aYW/HubJ3ToDMFxKSu
DolEqngP5uaxHuPduwQlLLvLnTKk5JqGaZtGkFe5CyPMZzhnQGCF/abSu2BROKteAHTmqYD+8jYx
5Jcj+YgX3Hze5rm64/t/kYkYCJ/7dTtUxRO+TC2yOzAAGEupw+cc8+qLLjWixiYCuX9w/n/PDb01
lgF/jsYaCGGtRjotGMugUeGhA0KKX0jtSevIGsYk1r/OF/jnGvdA0luuhlBuD0OrN1tSgUQ+ggD+
5MEyo1GSow5ww67jcnaTuto/xGYZykKwwWbU7W5ytNBWFtd6Bwl6ZJQ0igHkaaE1Rq98wTAbDJjQ
49VKARu6JlzZUv17e/kUEi9ISZUi3klXjxYG45NTC8ANR8cKsxRvlVQDADq3Gn+sywNPzRpFRDiq
StH+KtXWJzU8jrIObOxK8cbk2csZ1EMQ/ElkMt+HknBI1GGt4T0N/ToA6FKA/pqIldQHiMNROmGN
XwIfQKLpKzQqtpt53opbXMNTEeJ9oGN4+XBIbS1BLp8PQcFX+wa+x3/k6FTzU4nYPC7D3AYP07bL
NyiTto0+y4mMp+MuNOwNmk/aokBoO9t7Q+h6gGOq8RTtAmlC/GARzZ7qHtupgCpwO/XMAY7cFRt1
V1a/bYItoAmhizbdKBVRVDrYQje4J1ZhafMfAcKcPf3ZyEMyvTxEqh+ZUlS/2FIS4kk6435cmS++
Cbt6c99EksTACL9TvmSF1pwaWQDpaKqMw3y47lhiyYzrZEbcxKXtfv8RThi7UB0QE3ZQNfRw1w7G
Gcr6BF4VOfc++1m6nr46tI/HIGOW+4vr0qpmxSvxUq2KQwXgg4YMDMGXREEIBG+j8KimNfhDYaVM
ouGykrb9mYsW77xOIflZgGuxtOc4CAKX+SHRhyh9UAjU1OEBiWfKAF+XtsBDVmIw5fWjzWYA7IbV
cM6Vo0WOqlhL8jZ+q8y0VwdpAdCqx+PFCM4kyVxKs15UIGMVXJO9wGTOL9j9UjawlUAdb4/24L1G
vwvZn9zIM5KXJAod/WpahA1wO2SaEjcsFb+w+97iOLPO0zQ5MpRCvegDt5luJViFdr1YiwGR8Vha
LUhIEUN0/ZJ8Rs6ZpmDY9eFmPkY9U/CRStdhhi4zmxChjDZGCzcWrAQvwObetwX9Ow+AOpt5MBIP
Rha1DEfFSwPciDEeC+r+AOtLSBOVS6ofdIkRQ9YHHdXSZbN0Ffa90LWsQ+d2bHFqjJn7SBN8AdXB
neQuuLrdBKfQynIk8dzD9M2RqxO6grrD7SH6+s5quLRETV2zz+S66qlD7fc+sYroEtXufwcBK8pH
qweNzbcNCByseqGe5teZ21TdjB2H0Ci8qPjkzY/0d17n8R2jI4e7PlaoSGoqG6V5OlONpp2q3GiM
2/LST74jtbcvfaWDCdTDJTUumr9R6Wb6/yRDoVysMVGybPm9Tg/HHQ0AJ+6G2uQtRMob6hXu3IGZ
MB4KH5+0NkPVd9Y0RCUN8yHdjM2NK7vXat9My+ZdKYurfBKQ0UPNxDMeTuxVkpkBdrXJodL2Yhfm
FK6fYRX+/lppJOJOe0BZyb3DulKhqZ/naIG//UoG7NS/x+ZhuWA39ztf1CHnx79SjeMySaoLMKX9
D+YgBr04IcKKgDiziU7SbgYPIgZmsYgUinn2X3/GsnpBKDAzRLxFf7VogzFpK7Ah8ScYbgRWBe4W
FZaMoAKPcDf61/F8jHqoZhfyPydoOBw5zvnK2GTLhB7LAVvogWkwjRAreItXojyjIe/sH7H5l4zx
4IYiJ/sDtoumRw+EUuvtu2CyI51RjMoiAkdgmUu5ZHed9KF/zEQ5OogAc0ZmwqQH35NcNNbUVOEU
0sZB/dbJaKFXijxkQQqz563bwG/8yaQWeE19qbNj6+WtkX/YHdZWpJRNaYIWQVr+0AElXWkC98MM
L32uOYRwyhTcRWEKR1XmJq+A/cqCmUpAf68WRJN15oboAuLM7WSOHvAieYYqRgsuD0OxNWY4Rg8i
Hb+Qw8uF/TH4+6uBA89dKz8BmyBF5SD50L7qqz0tPkuRC3AHm77SrzCxo3rYDNzMLvXkpb9EG4+C
fPBRjzjvFtWfGleZZSwxyr2NMnLkFnpOOAZctM6+qz9Fntnt5U5W6nHyTLqnS8G3KY7LWMhpygRT
93jAmWT03einf2wx/+ZITVTAV4WhI3Ek8QtZJ6otAtDuLF7DtwjfBNYZH/TSjUxRTgCgihXn59ZX
Lk9rDB1Ti9R5vNBZRajJ3Wb3joTwN8ywNXkrfWjdNWDQ73G0cIFGmeAEG/JIqD/sI8uWD7zPnlP/
q/IxEESbA6AcnjeEyGKziMc1as7+QzDuLQMthDr6+4ewSa8xu/tu8aa8Z0sCzeyoiq6uOEFPmHAz
0Mr3/NiwoqPIkhQjL8pYmL8HUROqyse1jPq2/QJlCJzSQDdCNdR+kHs0N3SMnBQ06DK8g6iqjsMK
TJW4q4dBZvwIPFO0IccP2zP/ZFiYHn5fOBvZuXEWrFr1ySny8dE4AsdrdveONsA9TqCVF0gopnTB
hbNfvuIN2bCyJgdgKBFZ03Z+efc5o98B0loZ2aMCcTT39MiOEhlkJNWNEImBT67hEl19BcKdXSCi
TuvoD2INC7FDasNf2o0BQ8cdVyVlJ46UUzyv8xNZAMHwjsKfJZplt1N17sDWGHMEIfOFPjuu0Dip
lrQz9fHPd/1dRLsYfpCpHueoADrxrwmo4/T1ywPqRHzVKzuiIdpRjO0q2lYUFhZeZ+o/5a8tr1WM
u401MCDzQP3nqVk4GFoL6GLfIrc26rwaCBsnLmW+CEdVo9XlybbhCwHzdd9K+cl0ViCzoatBCS9W
zjQ+YCQUhSYgI9caCqvIK5QfiqpdsoKf04ahCV+CZ+8Ze2Ktp5PPxAcHTIEDgikRXsvw9ay4s9bN
xyYZ11POoY1QLEtUHULPlYlYC70pUWF+H5+tCbCy+NPs5MjAp+yR02wZ/tImptZNkTsHNNPnDypY
XKLHdZMdDlqgw68PvL5dCVIF9uB6SNdA4uMPn6bXb18D46QYkaDL8+nv+zCbn0FdPb6WwcKb3tCu
AXYStW5HSbpxTh185m+Xq1h+WD40zAmksR0UdAGrnQOvZNlJOy5TnHj8jqREbd2BZB7lOFZHdIsf
axn9uhbc5ka+W4FhdvxvdlkrSAEHx5kDGGZ6vMGPTaAxkbnTg9lsvDEcK994SUH9jsgOpiortF2h
2/cMvX49+Wa2pWonWeyUSU18oDtysgpJ5i8g4jXkG/kSGkGe0/omlHEs8JzKX2C8+/f1Fm7j4FeF
NnfTKEI2nTEOHKQ6qUCRtGZR9Xxz2GcCJsJcsyW3DW/26EqJFNf+uWbayRaJsLgZRMZNMtaXkMPj
0JxL3LP/ofn36C09VvsGpSQzO8cYePNg884igz2j224PS1i0sJGc4oxh4HabQh53GFAwiaqpfIQZ
zpqr337zbMtuo/M7+phVgeuG242VOHc/+/qsAtIIrQWi48BRmatsOsPFYkXqtOhZRvUpKBK9qxa3
+aC9v7WsDIPvbtti+qrHLdqTj4wOufQ6QKoqtaevsFdj1kl0Ozgaa7f3C7KIdV+OL6ndh1HMpv3f
EQA9EbqZYbDTi3BlSjmXdhoyYytNw8KHrCeTpo6SYTn2jpoZpilgetxmYwu/ZwpsjcUBzE0au+Jn
Q1Iwn1BlMUc+ivNb2yOzoI1vNEe2NnrvSQ50dd/4hMrMacS/5QGSfaR+fl0enYhBTmQfJWqj8qId
oXswm3okIw3ESaOW8y/1IX+GlV1OhVMhZeZ0RVXO1C0QYX5cfWDkkMvDVMJqVHch8EaFLX38FCCF
1bgpu+JhI8HkLWbhcRU2hwPQXfT73d2RjZ3qtNWHBXjodPKnB1omkvbP6LovmaTWhQUYA8zXaouB
WMm6H8N4dT31hSDJHqjqwxCFJmqCWBe3a3LvbO1SM5it1KcUCSRag47bAQuJMldrV2NQb7RoOd8T
EUU2kHynwscUP7XuB6W0v9EgwwS0djifhy2eM76gEIG59UovEaTuuW8QPbIG4OKz6JFh/1l17kBO
gV5UyUDcjv/QBZO7lX/3/uhG0ad1WUJrlEShPgslRf/IISEM3iy9nfYmmYV7qlb27704hN+hzCST
HMhrJtiumfRw9oYplh6MljWFWJtx/ipJka5ph6MtJrd8U2oc4qCWSSQmBDzjwgrOn6w8PSwPj/X4
yYXkoAH7odXG4FsZZ6yf6p3xQyNcFKSfD6xqJZPE9BGws4NmiLnuuoxorzzHiCIlnkUas3eUCvAe
SkoDrmuOpAc5W01/xkP+/CbC47HzuPiZI5sIi1EMiz/JLQMgyX4zn+LhdTvPD5GgXz+7TCfvs7gj
q6a9k0AJg55Bc+Uak+No7UqVj2kvdTdOvdnmZxzvRMTW3Sm0Ofsn/03JmomVeOfBga8aWP9wviEq
yuQ7DsQbGUvFHsyaVQ1WmNtJB/uKCeK7tONdRtxv8mCHHHl89XevVOlnLb82NC1ozewU5heee6B7
RxzwxvQlBQc3MmT74/ZtZAYemNz2EYmGtXiAFW/nSVrTVhR1ew/U8hfNfwFP1DKwqHrh0vzDE4QC
rVhxhHuAhwCuEBJcUNQFnb8Kb4MOv3hkijiBTd0/2x5IxiuAGq62lhk5Vltm5Qm7OQE0+QwRb2HP
uPIfw/1mXMni49Em2SLnUQHuLAI7hVCZImwIGlttTqWglZOi2IMLF3utH7iWe7MfpwUXwUTI1UoO
7C2nTqiTJ6DDbKbLAn0KCDwIVm0GHPGk17DAaVSjmuDq9LhCWrvpeliw13TdS8THIUBhJZmr1SaK
IfzbvjZLdJcoGQGqi8Nm0w1jUkU40m3kwtKr/U9rMq7/rX1RE4zwSTuCxH7cE84+nxZc/2BkiAKh
UeZvGVbT9Dg1UE3BmFp4sQGyhJYslmC8SJ6t03oo4J44BygM8jbFaFNSGOS6u0kn3jPqoK/CO+G6
Z0ykGuxJ7/mc+RxBDJqfZiraVsiGVhpAVGgfOe7VebYemts3EhK1aBUwWzmeyORI1MY10Jo0klYg
gFbOE6CD+b4FLqWag8WT48dXyXBPu00cCnts3TDY8cG9m5BwpcKBqk4ggtodWyqIhOWHgiYVRZgD
/zzLpo24LlBPZj0HZOavSuXrm84uSmX7IBbTbt1/9qJlD+bheXj0jW5Bs2LqTssEKb5SGfOCI/DY
EFfKmHURAEttmL6jb+vBQEUxJhmzGcz+9E9K22/sMA6jhRynGbyOnfitRElNbAViWvymjuyS3g9F
Z3A65BZQGSyUtuPzFguNWJfujhv5YHv93XatwfCzvKtUS3Y8oajsCiShktUcuLOFUoxQ0Yv3ebhJ
yxdYbYpqYUG8Nq6Xd1Jikok6QRceCtOkZmKo598m3h+xxsk1qrd+Owett3mmNWmdFb39LH355WVD
BWFWpi95x7BZ6ZCTACZRJ2I25ViLzGbAMXCElACZXaOLG4zA3P3FAyAskbLWsPXb55dsqLDY2HEn
LzwAlLSxLi822rdNERhy5GdoDFxw5LL4ImGPDMYgxhbrZ1X9/mY68IaV9NCqX5MbG4gepwOnsSfW
fPF9r1e7gqKqozHTqLjUJBxDFIrf06qt0JbSQiczpa36m6OsqW4z5bIggKHKak3duy3BsL+3LN8K
iINUxJQ1/DYL+dYlb5Ru8UrC7ZelDRHwEwkAUREWcckfgPZLRM54aRT97vG/iUnlVl6BNn1hojQp
o88vEndvP6XNepmQ9FSDDufmIc09IRwtG/DMcIBRCIMZDAtRd2OgpN9wcSFs5DmKOTt3NCRDsrlk
a0KqrCCV59ZEsL41rHqwjmnZT+dx1vrsyq4d2CDlHntHs6RhRjXy0/BCkkk8amTgSvyY0RIdDPam
e7LC0PkAJd9joFMxf2fdln0k1i49ivQwMCav6m0Nn0SJ0wSsR/WW5KvLwlgquwWzEcDCIe9CX41q
2MqPGCDwUv3IO/s21E2hzyEus37NSZQHRZVcc/iyC0kF5RhB6p6rWhmmIfbPbG7byLdZqzzA9ilX
OmDPIZWdrs1JSk43Wi8K8p2ddvRrLIfre/Mw9Vp52bTBYVMhsrExJqMhQWrxSWa/neLqaxpjwiFf
w/tqCfid14LGb4C2zis/a/1ZpJUjFnGlYjbCGilwkfwEUNP7kvEGQT8HMtuXc0ElFyxRC8UIA+lI
r5SteXCCY4xOlvuH8eCHzdpMmtjZu3OzAvaosKC+1JMoi4gE1aKul1TeYv91syXVHnlrk5DT2kY3
PxW70TGlmOoYXgPwvi86gzPp2zKW88nj0UyV0Lm1rAujxF+wXHXGTEoG3sCqBoIdOvGt7QlPFy63
M+LWV8658agwk1ayUNBAXD0gr0AxIfxv03BEcxP77ffBwH0bILlA18Au4bZRfoMnfW30ZTytGedq
lLkLp9xzX6fdPQNMY8ulHJkri1ZIQIFGXdl6zM3oXkl8cz+WHpKLtYnrRvl93KlJYCXrgyYSZxOu
b//5KdC2qim7+oQuTJNEAQTCdmtP1Jhgv9yuXW0cxK4VokkCJs+ORntrj1UYeqihye9W2QBE6rZc
FOYhL/2CVjboi+XcP1lAYphhe2rqFxbLvjhHsZ2nynNx1bZzczZel5uRqvTmClrCYXWOc2Am73Ke
koDSy91s2alYiEUCLJUgqJ4k7515xkzR+TQ0i8h3BhmowaZK0HRk693dwgsm0r5o3MqFo4F0nYed
fPjkUzReXw2lt75AxFWh7TOB9PIJ261PIXLbcWtSKpA89765gq8Gn+iNqlQYbX1S2GE1Gn5zdj9W
EsRgAR1y09lMfH2XSEMN69z5wlIXKsvoYicTFQ9T5fAw+q37gIeJ8nkFcZLQBxdPBMvgC4RF6H//
YudUeCuVzgojMOF5K70kK+qMP0eLOQjh5smYCtX28h67llLtxHMoBa4MFOC6EQv9xiXQOovwlyzw
7CX2C8+ILmuicjcNwsAQUkjr18GRGyunVrE3NgNBYbS/G0xv8Iplva33NJ1H+qfBzny9aZuseDE5
2zXy+odek6JHYtSVYF4K80bUrUHdRi0g26mmjP2p9F8tHQbxh5vB9A427j0r9vPgb4GxtXKekD40
wy+0avYfvmb00ZWzL19B1oqrCaau9/6oLDiB2OWfli2sMljAcVOqkElcoCZA9nvoggDVAvYAFQ1A
VnLVLr9in36iJvhSPi+Z/dY+phq5NPw4Rk22WaUhbgeVG76gDA4FOZBAxlDNKH0US+iYr2owN+pr
YM/dGox1DnSsPbtKM5M/RPh7OeqkzyGO3krtYFdKz6oh7L1qXLdELalvj0IUUZtnZX0iiTd5/51C
UtbgznMi0b5IEAwZwbb4jjBMw+s+FvAbfiT7AzG5OPHYHZz5HW2Gc21EgRrOSVl4g5TzZOaa2y6F
cH4Zuvuv1urmy7EgvevBkuk48iS/S92Pqe6re16eWe+lbRY5gyd0LtZD62HeHD6FFA5cYsG9/Aqi
7f+JWo42HigdCXDew/M6vC/yXmIIelFzaGoLwY8YthI3TXNR86uCzOhNSl/nL4b1tGf4WycPWGZk
D0uPWEGfamS+csFUjVnggKXYkFHO1QyimTOjj5+gfe+11T0TUP4hnfSMszx3lE2UI3bONvQZd6pE
ngPBvRoxj/6jMZR3lXGGWl7P0h2cDg8B32917bqEzsMFlPsONcKYogb7nDciKM3fFDpIlhEiDqt7
Us5eWvYkfb2dhSBNvtBfE2AQJzLZAvrTJiG//rV2OkfCCyWTQECGr49bHBODU1bF6vxpAYrVbrqd
gC6xbc9c/W/rQjJl3Htd6sifxDuAaGVBZyXmyxVa0yRohDFXWYTFtRBKc5e2yvWvOLiCfynX9Hfi
K36RqZqPtYiqJmIIW+NfnY0chmWP+h6z2noVImbxlYA/X15ri5OTyIsSYT1ZUW9+OMsR1fpnhj8F
36AHO81N7sjs65EjBLMofmG6bDLSJoV8twcaDbyCAbozyP8NgjHQL9qel/xB3V3s2YGB8n0UV7ct
VoEFGkUkKagXPwCIJuA8xt7C1ZqipC3Aobjn4oOXhuxGIyIbo3hGDjgvE5TTb61pQ8DaV9L7BiWF
s51ABwkymqI2rhOzsybJ4jqElISbzf3VeyAtRYolUFNyB2rLFRdhEL+Kam8JcVQ9QMrrH2/HapY5
dC1AhuHKPcTabOuTnAv6SHIuckwDziQzSIFOfKUXeYHKlczwiR5WG2+nhfSYsAO5vZA8qvKWG13b
NZPax+wxBqyJq8mvWOMEkijDU9A65qYuFFaKAzQzJbNnp6BalMntUin7ae5wOI9WMCpoGsSF9sbO
kAcyAD2JZ/jQ/IUG4Eei07xQKZstFMS7XDCBoS2AMdZLMP3M4GzLlmqmpx7EAwLye+9dMpOZKiVw
x/Orju57ARtyHBJhZftHHeIMRuMayf7K9/GCedQP+iznMLZxI7R2YVjZY1FkvHVn8EQ8t4ypvXo6
yjzQ9Mt+Ut65W8gsp/DIr1xfJkQy1osiVDEWM9qI2XfCnvQpsZ9dlbfdQvuLdeVoNMQkzP3WlX/3
fA4F8INYgGX5snATsnXlufKyMRroMWnI0XBj80UKYINq7DC/qM/DZyuRVBOgwm85kHGoM5syO1rz
4jpWG7YybjrymHJwKeDGo3JuzgK/umc2Flhnn7DcW07m8IaCWF+Z3KnKlJWwJd8QfSCnbJXLnEoW
lvc4+rObbHWiKs33ODxy+nXquItm1eewNF5+wPWhtn22RSi/wVYAd1y1w0KldERHFjJ0a29+S6O/
kBmPLx+MrlGtdppQHSHrSvVBsVZ7bgJaao2FDKUclr+0P51gxUdX2lx83RqlupbGrpa28pD/eO/d
AkZeuWPVprIvR3E6n3hZx0Ie0u1HW90zjP9a8ZeGXdzlNIPdVh2S//jnTEGPlkRjbJUu/2nP9YVH
+nbCIfP5tB7kNS4uA2xu3TAVLX+I7E6Sj4eIlkA9Qhe0H9/mbOx+06CwhE5K+a3xPm0wsrOeydDR
IOKHdz1lReB9OZoP6dosij0mm3BNrXexUzqSXImESTeCxFxAndVTkRphXMIZgdq0dwiN1z07oHZw
3OHTbPUF+ROUA5qz4jQGKL346kw+5wp/TqIAPGvEmMv5VNvHHHqr5bsRvZuv/wN+QpSvYLY0+jNj
1Rfm8BXvP+2TKAxVc5QGZ8tiE1YeedTekfhFTojlkGhD4gFGJcej+DAmYBFdVwR/DVPC1GPKWYSj
6gCKYhhFCRpgVl/gDsma6M8pq3TZFO6mCLGrerAnVcRqaQjqSlIohWyASyMPYt9gNi3kPWvyMI+s
jnDfNIlINZAVmUNJOtWSCBJY83RlTK6iWOu5v1yhYX4JiO9tL1sNuSUDkXKZngcpkEda8nYdVOa6
zn7pQCUpMAAp1V1tYCVErkgGImTX+ClTGrZMIqR4rtUPQuGHmU8PnH2/rENRfPX0ot2BHNBKWDSS
DxY5Y9h7lJHr+ecrlohuQCWn30vocvBhUvV4muyI7mqMfOh9zK+OfB62H0eP8y7bMduHSNMdyitd
1gUS+BURfGpfruMOWYeddvCvxK1pnTA5h3Lxjxk/x/mPS0s8Di8ph8typ7Uai2ipTULUgZbtoSLe
o7rOvBjWyi2Ua2I5myzZEn13tDgXsXrEGu6H05Od+09yOV7y0m1TZPFLnjhDNQ48h6224mHVdd6D
Fn6Ew4Uusq0GEG6x+WmLOEtRYc6ZdFT2Vy0e8LFF9YYqaa7AwdH3Q68bDW0O7dOzwhocx5nTZjGD
w/viYHTOrX26Czn3OF8ZqEJU6VWUMIjDCtss6Nwo0BQxVZVQkDj3cOr2o4hdG3Q31tza8jUFKsbk
xrHaQ1jWoaJuDFbu0+KFqx1XuEAuyU7ClU6FX2m+1RcvOKHGmRQXKykkSN0Vu4zhravRQorMvYXR
ftueskzPQp8ufSYrDlVrEsHtiytLj4w12RSyHqy3qQS30f/GkULoaiXeALjdw5IzU0JYakGdRSPk
LBqSWvh9QTyTTZhkdO8SAzvYDfkMuqBVIScJA6ZuTaXTzVHk6uRvoKTJNQA8YCTKnQ8Kmigi4FW+
mgq9aLjb6eVwmJ4g/T4jKIRTKhoGGsFoksIfDnco6xNp1Z7DqNeISdH3LnctPGzy5otbMtoaX9Si
XN2p+6Bcl+maZ98OYBg+wujeY3ARVfmidi2RxTIvVC7MhxFEKeOKeDwWFYI5hISyctNTJShjLTu8
Lk+O8oIBRFAPNuS/EkVnpQ78TwYnLbW1FGWQjkD96ZnkCj1ZFr9AvXy0SIeqSLGoulnYlxNk1DZy
nfso0VpERgwt+DCRLJtvo7639QtDEHgrL5e4QRJNv73XfWqo8mnh+PCJtWzPKsTN6WKPYLSl1LlA
vCf3byd3TzK0MvildC12ZUVvG21AYKRrtqRx1d0LIFXKkGg72Ujr9Jw9agC3fWfMAEup4xjk2g/t
Kk7vZdZ+VNoso6tWuBXzEFKbenlgXotHR951vY1rLc7E3CO7Pr29LoglJSRvXpcSnME2dT9Wyoa/
mlBPdoBO00VV/Rt490fA8b47lEwimDzoHDdQvQgkrOmaxeiWezC3v5HHN2ALhXEClyj6oKicEp6/
bgnH7e8JBMQS7ERF2F/z06uprjsDr0uy/xaW6JVjF/J6dnViRYGJpu5zGlX6d18b1dm9nTd98mQU
GeG1KxBe+COPLMyRtd6QD3KRYKhaVqlfXJVOMFKlPp9dugJEiJTW8xigm1mzXeg4lWXB/Zn+1TgG
i+rFw1N1QJN/G59sm7XAIHplfq787C0xjhSwHoHMrxT8M6gc1rabaWfP3HRIt/NE8zbf4ZPK4Odd
wKcLXX9BD+B8H6fOaGJxwTsL3ZJRd8EmxQFAPq7DDj/cFlzjQMAteuWw/NlxP09oOwYZbFkkZD9u
+7OIFjMqPOKSSl3y4C7dpT5+yCt9VkIxiITei00fxkZOKKDoYEvnoPNai5xEkeAHxWR1osDYlc6i
nT3K5AzGdkKPEWgPgFlx9yvr5vAdHVngV7K0hlSaBc7qMxLS9CH8YZhGQogg8al19TYxZGuOtDCy
72M8tyqh2xf992DRYtQX7M6JsuL5IS/PvcNocv8FM2adCjhKN8ABHsqCVPDfwOnfr4kDxEi5oUMN
xnr7SRfhfmuGPp9TbPFtyXgA8ocbZqac3Rpoam68ugeEWt234/yb5BDg7oOhVnioeyUbGXq/K7CL
su3SiWbki0PdjtRPT+MFqR21onEGsogv92Cw8tpCYzhUuYVABuvWz75SpIuH2BmnPZ4sI5M31JRg
kHu/x39f1Jjz37XFr6dR0wxpG29WylsmoTBhy7BznbJsOTx/vOJFt9lEyW939Ax25BUr7VC8oGSn
zrqAAi4gGJxFFVodR78dxtggkIihDL7LhQp8ovEvxu5ARn0rnuaUwrUFC6MMRDBUwnt6u5mzXyuN
uSHDITPY+DnSNJpksBuAbg3CkyA3YPehh6WCjZq3xqQUZ5t6ULuTtxdYq99/YucyScPYtsB4mOC6
WJG/OVt+0XBSS/Y8j80lidXNMKTNLXE5R+rwvFycdHQdlF/SbN3mSNJGv5gMx2pRHAiRHqfSH27s
+6XgKN9dukhzgWc4dnxXlWX9TfrlTJDN9/EcjtEc+ZNm0VRO2dqswH8u40rV74nlXv2jXHkLtHKH
zxLmELD47IrCY/cMHeJFxsnu5kkef8P4uuYBwNGwrPDO8X0lbPBHSlcKrzAPTpI8x/82oGJcTqZd
j47LWMZreHmlQX/I8vRzzYXEXWFPcIx8cK/FNZcecuBrVVzbxIvLn7AN9SKIdWy12+xmTmYwJ+Gy
+lGW2zcNZ/eseBdll8iR0S4VzxM9NP2bC02WNB1Nl6kN4fYuiRYM2oI6FLz0eYRfvahJlUPW2xO9
iYRUfPb3jDmfmk/1EYkbm4x8qn8z5f6vnpy+HkvH6RljhYEsFC1Ql6fBlPG1YHS6icSgoZMvkIDA
cjkEWSOZ1CpRWZcRyE5w1EPtvreQxPox43S/1dECFIwjujrqiPKMCT3fPSxDvCLzrSf8AXRpiGb8
LU9y9qOge6uBzaK2wx3M82HBibTXv3il7rO7nvFvpSJiUhHSigT1ZBMrr08L42LXgBw1vCem9E79
seli54deyNVtfll2AhVpAKxNuSW7IK+kvMDSEv/xAHivbPqwcwP3OKvmJKPEjbfYp2cl08cZRsm1
NZ//PBS2SYd+Lg2RMEzAuqkYrYS2PjXOtFf4Mfi7tY2O/abyfIEd2lBBewrDwfkK85zVOAYZACX7
rN0MYXR4x4/D24/NJ67zoh5jB0m26Mj/Czl0Y2c4LZIdvie8L20/jaFyD3tGz6M8S2MMRAdDgUXA
vhZr+eZkPB8sNz4c7mmneFg1lBmZYD+rHYHDiGA1Cqv1sEe/SB/iiu6rLAiVm+Q1BI7F+gIHdR57
iUKX4PxHQLN9PXzYOs+ne+kWOllJY0W+CLFuCd3fci2flzTzEJXVCiDir259vUQLmu/rrl8MfrZc
++pQBJSlkLQqgLAmFjWk4tdeIWwC39mqaXHa+aPmPrDQ4lX4XLIaHQqW0E2Pm9lWwhR1oWyWeac7
3YIuXVzpnMAHDFGFLqhAgQTMLn7nj5XWnf1Ra+foM9f3lKmJUVQLSlQB7ho3uBymgk4O07GZaG1j
/66rTRDb+RpMSjbdmKWTTJxqdvQ47a7aAP/YV5XdeHkVNPp9Qaqm/UcFYHK0O4xpcwiEG5FS0jbo
9Ludn4LAYn06LUekY9l/gYRzW3G6Vjzo/m/3vl1waVNhKtZIDrgur/Qbp6pp+atFC2MpPLJBv9FT
X551BE26t3QRkqdu0PB449AXsmGhX8Tj8Ti9RVv2pNirdnWKK3Vx3h+xrCCwjN9v9RMuIR0w7XZ6
eZOIZ8QmGasgulZ9srbEQXjIIL/KXGk8gatRvTueEtQ1TTSDOkSx8o0gjojHJVEt2Z/47mf2Foo9
XP7JGGTsAwGspFUDtl6M3c5oFBRi1ldEIRMGdFlj4fmPVDxOj0x73fqqrKeNIyYd6oXpFppazytN
JQT0A8Si7qUPHWFENPUkp9ZCGCZJAQy7uTVW8GiqZl7TWyT0Q7NwLNxLDiDRxnvxUl39lE3t5gsX
KrwJUlMvdjCB/lXDZ31eannRTMlm90owKa9dmcQH9GYXcR4TgYhUlYerL/WUY5vCUu1fZ5+RT22s
BK7T+o21WOyrGtM/q1ewMuyXUHibYn3Rq+x7HVer48B/3g8WqTNUZqAMd/+ST6tewXZrPX/XjYJl
4fRFNYaRqUhmEc0aOhGe+Lbloiuwn413dGTwQaix22jk8QmpD1wNpXzD11XlBVjH60pSQ2BlgfZj
d20eBn7RVyQ0ZfVf6aX/bJrVPldo7INdelbFUi/58THHztDif3F34y9ofOoB64CcTsah2Sagp9pZ
Lau01UZRZ8/cNnzleWxXxF8WXXRLxNPBJdvcZWbWYLm5BiP1r8mEQV3Ak9kaU3c5qb7nEQ3TgAel
qhnXilTEwLWRYcWqO/hqNoF+6Wob/NiT/xxvP1LIY9M/0azOV9+kPuANmTgq6bbRAWL5Mg9kaJwo
NTb3zntJgLtvR1laa7amhdbjoDsxO6wdg3q11FMxjN51j03LVPoqAi4CBgUG3rpNALkrb5123iXL
HGhl0SfLe1bRYOzI33Fa3l2dnXDSQMGL0rcsEl8fQYtU8Yk4hklKr4aK9ltiwOWgKZLTUGPTUkxr
n0Xac4ovMbmEKgLg/UDKMoUKz5Cyt87CJuD4yPidVmcE41pk1d5Kqf8ouxnBF1vT5dsi1JxoQPfF
0enOnDi/3lYn8kCgjy4rHeYVnJRzFkoxlQwFZAvb0OJEUxITsG/jxjq3A0tu3pyf7GHRQ07iJThO
MMhdnWayq3f808F6f/yljjxPGoKA72BTVyh9/uSD94XT99AQqd/9z1Z8roLAS4Pwg4WQDvcHn9cw
kPgQlOQIVZF3eo9S7yFuvVhnkJLg0f0rHJAi5gxbs6qFEDM9EJEnWhbhoohCJWOwFzy8jkMchTCf
2KAIFTGpImySK8aZpDs0PoHOTGjJ8g1mYLuWCT0B+pktq2enWzN43LT5ejIkMYVsdWwmli4kJvb6
zdIs3NPPScshYA37GHV7ZT4NtIg1c7lOHDC9y/UjTKfM3cUFvqn0XEljoxVCZmM/Egtz1l88Ub9h
Q7pQPYxp+Bty0xEoRGcFFQ+uaSla81yfb280qjlvcp/2o5pQior6XZSxDLasGPS88sT6dsyNJbIx
LI/ZXEwClJRFJFcKAok/4u7VZCJO+U08WjW0kHzoaf+YYtcK4GLMsXbzn4InpZeIkLLMmpWXPA6o
vmftidTTUdC7+vRnXcflrg76RCVX3lXO65lwmQaCqmIf7BMV+QHr+7rkg+EqAW/hiabIeleBKnOn
0fVp6RrYwLg5QCFllKsuUKJsD9cJQOaICnlvMSWcrVEuGBWc2aOACoDN3PrHgH3x8D65gpQaPmwq
dw2lcXZuhxUFqb3mUTTykKth7BlwciB8FnMbdqyeRUOMZGMZtFjLV8nNEdiUE33te4gp8pEW8R/O
ZPpYqa5t9HaTxpLvlLyivnofPo9ccp8NjDvLHki8MBFU8f9+hPqk7rhNozJ0R4JcsBWyOtPPuqYp
F/8NFGkWS2E0VUYE5S6eYlcAwtekjyYa5Xaa886ByEBRqux3buCYFSZHMVn7N0fU4E26bkSkWmuJ
lMdmFke02LRMhtXm9sD3OXdhKjOtiyRL4JqUA9hftYhUeGC8pNn7+FgzDpmfoq7ih0UAy8McdAvZ
h7T240zTgdj0qB8ncspsFtrjvoMxe8UBSS/XbBq0IncuaV3o4M3sSLR1hzECQME+fnA40+rbKu8w
aCsIJhjG+5R0600j8HcO1HiBOShwjbcFuPZ+gN/MjBj7dP2YdfrKUUuczxIrLQyQCHEYgoPaAS8c
Ah2g5Vd4t4IQcPASk2Zo3cbuDBHDOBIKm8lCj/27VmxkY0w5i57dFOkePsj2Y52M7uHqRryMjf/A
KeoAavLxbvQmJ1lY7CFnRUz0JgP8j6Qqr57rrDX73cLdZ04ngtYRKcngMN20hA0hLzK7eHYk18ob
if+W0rYxIpcwB+gfD9t3EmLzUpN/rhgXSvKyV46Jh5XIq82eneLxSfs1vKAcnuQWixOvYEutS6bI
KQh2eLxzgXmPg4ardmmWYaDdAZ0m0CcJFsBdHpH+4i/H5anvd3WIw6zcMcZ91KD4GKbH+TTI76yt
cc5mufO4xafSMjrYWUg8wRsuNDD0cu2DmqCMnNrt+WOZvRu6e2IP2LR3AhQGli1vFno/K2A37mBS
WSO1FnaiPppgZ3ieT0zyoW058DIvt/eNEUl8DPrl25xSHfG6YNmrJb41geWKDdnH3tiUfj7F5Oxt
IZ88ukwCWhey7GSysx3GSlSoUD5k6+O2mO0j/EfFwJUDLvaBH7c71jOlfFvimYNokFBvpYTDbjeg
X74FhKrwyAj0mVgmvdZJj9hS1+F8NOtMthyefDM9v0fhpADi/MOCu0Y0KKeBEF0N4iHGRKDortA3
g7EQ47Aa72jG3sFP83TADkCj32labx9+DoX7wNWu/yaPR6pUXF2oxihpD6Km+FLOvALNu/eJCPtv
qb4WtDcfFTMBdPjZS5563tckIIjumPEs3oWiFQrqBMWnOc+kQ73pTCsR7CGYsSiBidMkywhIpycW
KK6yPl6MeOIZzXIbph5uGjbvZ5UNFWMqvyhTHbgFmLJV0nG8Sjy9g38vBI5m+cBB8DZJJlXe2Thg
GcDBkBsIfHD6PGdt+yYiya5eSKhgK3pWnYveyGUs1RD67BPvfXniEYNn+YzLxD7c4gYS0fo8xSyw
XMJWb51yJjOat+6517zPUi/ehJ/s9fAQZ3LYKNyCDiljRNi9rZBMDox0H5kZHfthm5+UX/Po0OdO
Urf2ohFTVy8PTicuZTTtH8z9NNDbc6zTuTXIifUkPmJH9exnwWwrRtrWzFW+ZHy/vfzG8xhOr7pz
/zWA1Oo5SGJWxv/uUn1hQN13ZV2RLFMAw3RvG02yZl4gXbiPWGWS8Ef/s2r3rjpGxWh6OFgzHgoi
473RdHdrYQfi7WroCpuvnNtoCLfe/Fw86w9Ket8dC4NVd83x8BbbikpJ0BU1DRZt1YGSwq6/hCce
htuU1ErKY8jRJjZNC7afostFr09MhapSD6N1mU8zD2tiFIEEOsj9KdUvYH8jyF/yq/iVSU4+hscC
KDN+s8jgxYpLvIwSpZEe5SpNza3BpYhON8Ga/QBp/SxKq2jndh0fVtqc5OvLQMFWlta4K3cRGJOz
h6JBlDGPbcqyQXuFQ9wPcO+4RGoJXSntuTaY8RTFvrpHUwham3dmN2dOZtrRn6k8EeZMFPkJgpsx
xISSlWVjohFYRwg339umgxyeWGGJvNG5xmPu3nmVLj+LPDcPJHu3/1Ue3V2n6jp1viIEWRxsnbVd
OyBcnXl4rX0wjlG1671FMp7Ux8Hqlw+IyqdoiQ+mB2jB+EWZK2oDJLFIumC3vuBzUpCte5E/2HG7
tv/F5nSI0q8/FYGBMsDt+QBsqNO7kJhdYF06IKeYnFtO6XGKn8H6mdK/F8PakTBNUg6Y7f17TuCR
XNI+3Xm6J74d5xDxrPZEhDh0G7B3mkfbyFu67L16crAOyl3b8yWJfjdIbCm/RSG+EnrEOVnNPNdf
rxMtEvFLAePa13Ga+zM0FNbmL4wZSYPwBzyW1lExR8hguNMJsMvScRFJxN6fJakuRLZatqZHrXfe
/fYxHG0wO3jn2XsItpuwlXHNEun9dB22/IUHdi0saxBCukq96uK6pYSBWh0Qml0CrO4pMZDF0pNQ
Mxi3QqqCgFl/YjgAT0RTTxvJIMqMjF1ITO24FCeUHAVj94n/ScOv4rK/2iMyNvW2ae9IQVd13VOA
i2Rd+PKbbrwU5+OU9SFjDa36e+7cXVjm6gJ64fh0vRwiEtMjHPSrpLfTx02xdX20lZ75L/Wb6pOW
krwQ2d516S1v/MULNibzjQ7tTlpBrpb4AJSJGMdxual7myq+OVJo1huBWDgWmWS1b+8jd2oY5zAe
iDeJSH2fwc9XokgdMwVe92wS+LsZeC3ajxSlp4pVXU8OgyGX94xmaNl2AEaAztsSYjPT3ieUvwnz
7P9Kci+BxCGwcJKq+qWvNVzEADdBYv/7UJANU2PRYGO9+OLKQ3VHbwxiRpH/bqkgrPScOoN2hQFS
pb+dSX22raTxwJeQyDrDgyexGWRomdHxi15LKHvQoAoSzDyECmC0PZgeFqd0lQEN4wq5eKVMhpxe
iizjrdirHdetcBsBzYlBKoaCAgPAV3xIZ3Aa4BQiZBaVmHnQKlPbzPKnVepSt5PHY9t9yWz76xcT
9UqnyQnDT6BYhCDXZLM8xugYPNOAybFS4NgMzksVHRbZOliAuTtaWCbeYoCIsnncyQdAx3Hrr36k
12/X1VWP9hyCxsB44ADNUC0gGTIBFuX78XJM0JmiMGuGWcTnquCMfazVv/9acNtjMg01vL5LHAIq
mBDWCeXsv7jzvCjDk/fg86ltAe3QUXRgXE80UUWYg3NBAv4qWDKeAEEzaDNdUVqTvoC4I5ysF7rJ
EzTS3F7JPZFtL0PCk7AlZ/qWJNIxl9XM6pyDx6+D8eY0h7DNJNIyFHVDoOuGaUWu0cuzppmJ6rnZ
/ppbfEAWyJN0POvcMVBNpNywZe1WqX7xXXPHPHp37r/ginIIALo4/uA+2ifPzeePWPaCm8eL2iOl
0LOTuBRVyE3SapoLPChiiXiM6K/h0xDI8Erqqkj0ew7vQuLwDCUvW/rHwzMgCVaTUU56LOmybX/K
BDht5J/i/LNuVqstkV7EsX9nV50wO9PPDl1YiB3HMZXvQfGYAIem7ZBGTq1hLckcNIfDCZtSsieT
KjvEJmN0DRs7zXbFBT4wclLCHtxIuvrDnYYv83Tg38JqUlzpSWdBodZf313yjE5nuUNN+7iUe7Po
4illeyqlF4cP1bCvuxfkYFJ1GLKnpJiIFpiEXQrfCzoDO/p4ADFWe2A0jhVpQCsUF/xRxen9O2ce
arsibhx47UaLcmOISKoOPxtmPrFtdvvdzbQtiIXUu68oOSSWEPnOToAlnLV8qNV3Q2e1vTrl9piV
KOlyAkUUl6T+hppr0MWCCJ/hX6gNILinh+WmDrg7CwNPyXhuJyMgz8i7fYpT6CAkbdZx0aUQwx5v
Pn4/Lfcq0Ko4IyxLMJLtssaKm/aLCfZixZ1pjMi6DVe7ekdxO20FBAApnTnOihmY2Fg52cYyU7qU
pXjQ0ldNb4obM9v6oGov3Repck6l9zteM+CvJrUWCS5oLy+J2Ewtjb2muIwE1kpW5/hYhFdOtbFz
669brOC9H/+/L0UFx7KGMnKMxmrS/PgFF0A2ge5Ts4rCkkBIIXmJUB8v+ifF/MKee+sXuh6Jbu1I
hXd2r8kGBn0U3NInKiJd3Tuo96ZdWSTWNqCdl1KSRztT/HjGQBfXKsB1qcIve/gPTJ5rktPDpuhP
KwmwzikPEYsHjUAtJ7Yp9kT5Iyzh583piw3Dt0fKI7NasZyuqdHJmGg2j9ATnsR4Wto7J+SOg5FC
asbZJNLIGPgHG6uyev+CusXbFHKYmPPNbhZrkb3ePB/GmtgDgt9yfmmk6pt3SwNafkN361egkdYm
aSqUyUDwuQoCuS4KllsAeKt8UDy5O2qGv0matILEgMXs7tZ7TCjZI6uBhM+3p50l5RVHAOWvjhSz
AsYCXglUYftX6gG5pw0vs1Lqu+2C/Q6FZHB6zAlvE3GXI5O0MVZTkTq0jW3clKenAu/UA3i2g/z6
Y6AEHmlS36/lmBeMHazVygY1SXDFs4ui4HBuI0e54NzPCfWXwfRVD+fU2nNPJw43824zFi/tLKYq
sznT50wuyntHWNscJlnJcwTcwyuLjzUhD1hY5TUjouqHbO3WexFzDeBRRz77NnvMp9hTfma6img6
MgFQZKYSRkrqWjXL2dIM/rOeM+UKBmvZKBeAglE4ykvP+bZ0jSwywsTq1vbAs92oO0fWbB8B6r8g
KujMyqVJz29LTl0J68uqZj3b8Nq4h2DTrU23yFEq9Mhp82VA4KkRuGv07KRK+vOFcxcQLhMU8NL9
jaYbErptAa9AujiAdxBFDb/AevAEG5JB5w3KBOwTEDcPRTQslFhnO9aUnV2pMxGUfz6yKNiPqHYI
SMKlPcHAQ//EAz1WIchfVfXdw+AxbY8CJFZheFOXvh1Q1QhChGKo6DiMg2ASODFyeBPddiDpRUbk
+FtJN3ghyzoYhplsXYS5JnHWwBf+4d/CZ7eVj2DVJGyJHc7haiybutlOEiWqrLqlSZnYBUpmHXE3
LlH/WjxqJK8mkPpFFQ8jiP0KU5HgGQD1JhUwK7FTV2es5jdWCYoo054H4at5yA1XSYOBh14sphTP
4zEA6D7dihKQLKfvr4NuzD77JHBy4gK2i1GinK8CQ/k7Ud/NzJLsIqHuUc4+Z+8r2PgneeK8Cg92
Jn1LfTZHnIxdc+OaONG+Uo8rp0n4tVM0WsVtE4XkX4QRJKEnZpWZYQdgpbUqdgDC0XLLVfVQBnRY
8MT834IiQkmuI/xnrkBuA+Z8Sig7iM5P6ixvKwFGB/XX5TW1XaHewlf9fRTmuEUMQutUKruKJVjS
5fjxVttIt51srFfF+YIzoq5yzlaJCixtWY29E5FK2ACn6KVnKznqxD+y8O1Jke+GeYGlwwqU94RD
u9yjPPi2Fz5GaxYVjXyYBpdyTDX2sy0YoWVGtO7z/Itn2SYsSMMot6tWBrTDd/p+Ww4UdVzL20aE
CblNUHqS6fJTYkyqkthKsWurSY2ZM1it33nj/1dEhweHxHBHK7ge/Ca7PfhYrwUYL4B++hmOWeSC
3UkohwtI2B8Dpm9Rv3MgXrgzV2FIjXtbiOIM5XN3JqrMbBXsju/B9epNs8cF3IanPcwAWuqsM5g5
wecuT77wB50HMEu+3OgK8TYaKCsPBFerm8QY3OHZ9ZDZtMRT4F5pLzbfAsHpXPpLv8fXkOV/l3/p
pmmbrsRwj4WNsSu374zuTZJZ1DEGjVdcqZXokTkWhB/mAqr68F5kRPQO13dIdAZ0hoDLUrKfwnUR
XJqcLYB3nJ8JetDTLRwl+EYK+7eFh61cHMKtKhvxZ664GPnoABZnYhlgKvxLxwV7JslCup/RaPdN
1jcyMLO+qD+OTAbJlKqoKrxfzIf8ZB8SNJ76pcF+n/5KRSMa2bzDCo2Tb7+7+jMo7XinjNzqQ/Yi
Ttz6Y/TXj2If6opVGQzSWLZAeTkEkRHIr9ej+cXgvlbG+D7kxI21Xp9NROtsNuaDPjYCvMe6fPci
iNhTq0fCSUkYU1P3JxL2BZ3AEDr2M6IdntFXJFvwJ9HJhO5BF3cvpB1Ig2O1WDeZ4K9YlIYQ5zCx
hbOg0zFgj3M7P5WssCo9KUmFPGED6fnb8PN4C2FrCq630sZYmAG6A5ZzkR/o3IMEz+iYNOtHOvF0
N6DM/aQTZ6peaY9FISFw4WsASql7I63KsWve+U5Yu3EgDx8qFItcXLQDULQe1bByxm/2B7aOeGJ2
SgqWIVxMDMw2VyaKN7d89SGIOiMfauwSIlG2ZIXjLg5+C95ebfb049IUnl9CJg4D1/ahCDxYAveD
BfSFn0XXu/EXE/6e3YOgiE4IG7tVyC2/G8X5hONF3P8nazLLjC6EgnglrE/5BPPptHxqy6+LjOvS
lm7uhUsBPv/5kJz9covuv1QHeeSNy1eYHHIvRhFsh/3brt/RNW3tB419pFyFA6DBy+r9HaJ3you0
y++/WerbaSLc+WVTy/IXdZ84YW4/RPLBk48/1mS+hFd2ZU06G9SKAW423SMvw3qILvYdLTPaQhHb
dgHnLhOf1pTDYyAh5kNWxgEAPIrUtiy0qPRNJfecHAqP8cJC18qqmqfCZCCeIuasUj2nBwdhr86j
i3v750NsgnR3n4TYFdTfR5OFNuPrKqhVPeEVQ5KYMqw3IAJtz4QryFOkep6OdGyirrXwxx4DHFf7
4UfPexjSrsu3R5IuQxumne0QYPB6O9gxl9hZA7XignjsaxlaKA2et2dBW5vWMzw9Ygb2SDIHhm6X
HhBuK+ugBGkhMTaAYWOm52qckSAxNtzmueAdYl8AKeB9DSQ9x6WWrl2gr/+UoXpZzWPcp/opC0td
RliIBPprfnpLjqFdwlIfhsxho1ZVzq3rEV8fhDdJuqsDe57+3siuc7yzBYisARE4OQEetFfYc7qk
LNEYGR30M9CT7a4GQdmkqQICGQM9e9+p9filnI1EQQkMUnUqlIRfqLw4Dsj891HYzMD62tSLzFHa
qzbIUkj8ttw5xZ58W4o6pzap8qfHb44vXJR1WZmLMbzHaK7wJxxXEQNY9NJP9Ct8yWOP3PNl46mD
ArvajNpFJWN3/k50mZGOrT22KjF/To7A7eKGySdGaPG+cllkrYdkFbU2d/3d5JY9vmk8qCRnepBt
nSdscE5XYNfweklsKQWuqWwEl1/o2mhxZOvsOoRysxZki++eaJZixZHuO5qVP/hEzntePAzAm42n
xCXtMRuWgeY18l55kWRtxhAskwh0AnsvrLhIDoFxf8RzHarM1PHC2HrQH/acRgvS8i7WA43dMtgH
K5PaMEmG6AuggdmFU/hClpIc6a2Zjuv0cqUG31DOa1Cbk8kU24mt5dzr/23fI9jACqvidBVHePI9
wOOHPm5gvDgM+rF1MjFgrHFjk3YkWT6BMdI2pAQ3y1yqVSwPgsAFteF1EYrE8aAUnHXdlLmZ6qJI
aKtBFIfykmyfyk9/4lK7vG7W9ADHSmwBOCSZ+JF9u1XQVCV+bEPHXL7bweTvl4REkzyuJS/rQZKe
kRNtZNLg4Qe9vdVrz6QEv+pnRTPUTDJ0byXwvTQIq8vL3BSf7ULMpWJuazz8WF58tKqE0Ac6Z3BJ
LiOAIN9fEjrroZd2CeN/b/EGsKaFO5X88plG5ooKsC9goz8ySONdeUhps2ANkVi1MLfO8E8fiFDy
DjyNJIfY7gIz8GIOWbYyGfBCjbacpwCc3oudl59chh/NODj0T1MkhoUeUjszN4xbU6x7NjbSDQeC
6+bilmtHXzhmcQPIZrqrqoA2jVauhrZGyNUaL1EGPuz7uJFGmdjuwZCoFPiX61rYtDoNIj96ODbQ
KRZ8XvT1iqkCMD9wQQxUewOYHjqszj7Pebsic2i3Ts7uj0ACuID4Tf/JF7wRhZg8fjnHgsFX3dY8
R37JWhJlj3aOjHZ5tIRJBa4v3mpZ0zNNmuM6+caSHItKGiGX64zTTt5DGTBLxQV/pVO78cK0ITlO
HbDfYjWaQ9VYSODUYsMS/wO/T7Vqk1VT36/VZ7ZKPqWACcB/ICYnsvO4BkyqHCy5FusRbCVoMxdT
xv5aSTy9cFHfpFykB3pII1VEaLDUrzKqSehLoR3q1GodVI3mqNYUrkyJiot12x/h70p6FeuK/ePQ
fq3dQmn09dwF6Q4tMWxX6feTuR8SZOkXvq0b4b4aXHTchLF8yfcBlpK5VeljCIu3cwV8STbJDraw
ZuW/NQw4a1hn4ON3iuC0uME+sL9KujUWZtZO6FIX7pDvDv6N7AKT9Fo0jlf58dR3Bsm4fbtgVs4V
SnSy2UCZrhS4GhRynB5kOQYy9yBRWjTH1fBQwoiGYHFgbfaeHkEjBAmLC6jMrc0SBFfQMT/HOtcY
eUzEPNLVOslkRHFpXe+PJK3hdIGooC8sAzPRJFk1WyEOGGBOD971WB4HAwIkbLhMkueWnycl8Fu3
g85cPFp0zQ/878PioLSdQB3H1ZVivIsTUjab0tj9wYF66lpeA/D+ywFOBP9cDWWVLu+cfI54NVWU
cdMDmaRNTznx9Hd0ygJf8i3lQ+8QnANeinifzrP/x9fZ25x9LzYs1nUXt5lJYYiMhfi+xmus8qGf
qYtJfUaQ3xVv+Y/wgf6BRX9yQiv+M/x0CDUofLu87kBxDWw5iKvivlCRHuM+KQfhdISULjPWb5Q0
aF4vwMbkIHQqNeAqH3c1DwEYVo7i8vBq3NGeFYbnQ3My0wRP2nhlMXl1gsfk0XhLJvKgOgoRbYWe
d+d8b0Qn2DNoDB2GonulicwSLEdqIDcs7oTvoLrLKFHYZWFR/nu4GTDHhoPtbir+Z7osqopHK5GI
EWS1JJT4mkV07pD1EUH//ghN9LND2nD4IlLzETfsAXG9xlly5ny/KpOOo8Uk4iRcAcYC9H51Mnc2
JXhf5AIKOt6oJxnZdhMGwQol1Mmpl4NBlVYlpLACh5bmY1IroH0Z+EASdo4udVCR1yBG8cWPzmfg
1wiDcKxgUuAlkqUraiOFENH2N+Ut2BStY5Cyn1GjkcG7g34/EW0iOg0pM7k7WpbKLFX/DQd6R27A
Xa0+dkTW0FBggpSkmHFK/nz6PbxSlmbcwRdpawGpSGDOUZ1ULAHyHVag2fd5TpfmBcgNwjeAs2L7
n9JKVoMOk5DQ0WSs66zHZ7g5ui7sBcrAP/Ux1SD36R0z58R2xeMm8wW8wJa6cfkJJAleuBSXLPcJ
bW+XkcjEe4rVHj14Ez61zn9CrhasFSxYatkqj5EuGrrdkKD4/ihKBv58sjGQzAloa8pnWDOw8O/c
mveOsyfkSrZ6PBrxgaTz0BJJKYLLk+kqEVaWCouzMiikV4bmOU8ogE759jx1FJx2mDOV68/uCOnV
7SsCSDsMnAgoKgBY+72lUARVtUJabw80LVRupFAqGD1evFznXo5ru5KLCiyL2ek7Aa8fJnERIJnk
1SMYh9csLdLF4V5IbgQgBt0d+JqNhF6s/GG6Xm1SG2QkL7nke9v9p4DsN9RlM9vWMVoSV5/fPoCG
T1404uOiaINOIoVgBG7f1SSZFURioyVNCcTPnSWxdbrysQoe8QN+/V4AwIAIQHL+1sRmSK1ip1z0
EiXDwnnhP/iYJwdUPXkvsm1HvwQf92k53Y728ThPAko9hiKjROBrLdHrjj0kbIm6WOHKke6lTplr
2UgapeEE90wua1r0KymebyfECUB0KhNxUzajwNxPu2E/kZjGxJcbw7SFtWVLPciZVaBccGqjfBfL
yQLPhlcMgHuq0L4B5nqzdwWbFn1V2KiDLFgvQHnlk+R3i6GPcKQoyMhq7RvKC8UIfZpHXlA2g/ku
vVzztaecor3qGDpQwwUji+/Ni69Ql1pV2Jiwq2OwyZNWUhyZiVSL7T9IsVUrcBVTEmnNTPM9nJ80
M3eSCI0FNr58LvvRN324pXNi3XMXFlppitjYuXX7UcjOgucR9eJN1htmAbslW20MYLqZDV2NDe4h
eaQXZXiZFPYjSK2P2mYt5zf/7veTimdpSc5WwoT36wCYmqKSXY+DK6hfU3imUgFpE/Sa8KTQsz6g
0t5eckZfTqwl8mqa5x4X8odTJzk3jfF0rWgY1+M9mqCRZXuewd1Jb1+OrKhhOc6d+q+W25JuSH1e
3nRB4arseRu33yQNu527ZqbZPGTOfkSHVsaue4scOCBbKU9cdrkgMIjDdrsQllNwFs7dGpe5domW
JY7kXF0bIfWZdPgDdPQxoknzalF52q28GmWGPtZueexw850UNMtEvt0ZYPoJQJj1kjzGAk4bgjtO
yFRi7ENmfwLaNFfLqVuytcccSdNnV59l1/Bt3EJBZud17QiQQ9SJPn4o+PU+gqjooOCJmvxbCgDD
SK8l/M1QkzzjWSSquqvu0PRYi0emjjmxTBotuMhHeQ7GZbRPq7Y5vX+LYvUvzYLs0DjpDFgXnk3P
rLqR6jr8xX1nF9ejBqr+qObVjKGFsz+xPCy9lFhucyM6qjZRrUAb6ZjvGzfIFkKQCZPpwDAsNrTH
p6J0r80AxA0MouBBFZfWPRyuuFdGs8d3BCsgciurt1FGyVdHw0Mt4wol4r3K8PhVrK3xg4RyS6Zj
4s/NPYV/WlmWTblfYwpY6mMyiKznVyqlyPoqVFC4g5woiAIUXxsw4cQt9v0hoxitQofDFCc1xZdx
fFdpOc+LRsH94U8Vk+T/e/NABMSzVVRI7jh7s44i3JI9LSEsAmUqvTlPgrKoa/ARBPqe4R4llQjD
EDlXvYsfIdgcjkdjoi741GbPFyDi1gOur3KTQcusju/hpwRgeRltk4tqofjFw8orgLDCu4GMu6Wm
JMkPqqTXGeLd658LNPQ7/lWbPt0mwoQpZWSYwT4wgl4d8CAFJ09Asoi+suGA2s0C660oL5IRl/FV
q1l06BwuohPk52nFuaYget2M8AEu7juvZnGV47a7ANTyNTFPsBiWWZ9lAxjwuSck4fxOkxk1v+lU
97feKCW5Xno6gPG9XBaqPwvYq6mB+cXbUZnexO6ZDnU5Ez0oI8ehRonMwluwIA/cJF1G6SatQO+P
GWNBKGRB/g7sGZUvQQjW7g6BMhzL1wvNShYmHAGfaccF0QPgML5vNiiMAKExOOIVdt05mjV3I5Yu
PtXCCYgQOfGpAZtYVNE4EHg/lgai165RX5EXY9UAT5H4Gcx3y0nptKshvMySxglG+h0+P6otcIjE
5nF0Y0G4CkXNR0tsi9aL1xj3w0UjDqDZZqi/fsg3g2TiDXQsFaGCEkN9rFzQNtPdyWh6E5KWytY1
ra+M11OYisKwOL0uI65X357kt1VcDwgAAWSOHSPffTaOG692inpmRtGir65mMsvFrIGiDJb8I65k
DU4kK5e9cbKJkLrHuSc/p5zYa8TVh5oR/ILhct91Y73QSNg6xakBdgfUdNwJU7fXyz68IBugFSmC
iumWcQd7YfNCDnDQhyS1qFB/FddIX/KJ0usyydAC5STEbuu5oylyIK8J+w698Dd8kk4/6hLttatd
WOReNFkcDlwyfnHyc3klQcnzn4Rqpn4FQ+U6jFyFzfWfcejk/ZlJHWdf2PK1mWRZJfQY0uueWjh5
wkk549AREW6ofNG9CxCkntsAn4KmR2U0PwaBoOgRXo/F+/MpaqjFURFwi5zyb2B0kNvprVPDxsYD
WkgpvFmpNGFUy7GL0Lds0qnpTgCBm/raur0NL6vAuaZpLypqoYxEh77Q5WdgsLMeoJViuSzAAPbs
hnvoz6CgE/WUknfcJ44AlCKCB4KRZATxd8zvRgnHP5CvVGhNVrDuARr95RyZgwIIhlY1baW4oAdW
WdEB4ZmXVA/nyr8Ab0TMZM5c3s2yRp7J8LmmO/7WwbCjPwHTvCDrwz0M+5X+aZEtZW/vqaBrn7j8
Df3J1kScPnePARFdZMfMEpizZ0CROa/jKFa2/Eb8Fg58L0d2IMylWcVHBM871B7607VbcbIPsXa0
Gm8AAJh/nDkdbs+JG/U9ete6psbLEScCVrwZnHi3+KhQ/198LW3sgCmVtR/TqVPxbyXtxJF+MiSi
hyGKlh0tGViGXZhtfVxPG3OkH1hnxgfOZAmR4mAQ9jklXcVL3/6DTc24s1E547hXOelekdA1Lu1S
w/UJJZeYeY8MBscV5/l456yPlFoRbKytRXtu03d1k8Mh3HnIvCPfn2KBgJ+CdudLkMs871zDJy+Q
VzeejEF/EcRX0Y0qdVxIspYgNCAwVPWVizF9GnQUtJ7V8U07c9n1y1CFnmvVJCboCLz8QLGGSzYE
OAxUd6nTtGfx+w0bOviQ2uDeemyWwx3AQhiogepTUf1eDCdGBEXFTjdwKtMZByioz4Fxb2SfANlv
WPthXrCsTqmx4Hh8cXQ7R7CdSbAt9Ly8zYZIVTwYqcut51ZWPSYr1vu9zdBzw2uipChB6fyVWiOE
uEpGucccsatYJpuygYeTJ5TXv+XwOx+TWaha4qG8tHlpbPVeeUxKM0xPe2sAz56dyBAu3iofaXwc
rWzNJ66UAwBXGfLpFEUp8QDW6IQT6A3wQnSfr8UcunSTXt0tQ8uMai/xqxUlWrERxX9HDabirqJm
s/0f9oAQM8LWzL5Tkl4b5acCf9q/1Ai5XQsuXWRBSYPujJykoW1jH/5z6JiScwnglyXbJ3z7pVme
sflPnfY0vgTVJArBiZMGdms8D+CuNba62F1Ry77Dw6qX6pQuV7892SuderATYSyDVC2CdxDv8f7W
Oa9bNuoEHggiCwf3A8euN235xpg5kYwFPxgbYqvCNY8mfN+9xPGTbTpFhr6iRatdsluI4n4ssRhL
6BGZ3JtT3vkPDVhPGgHQVF+md9/jzY2ow6H9NmRxhQjIo0iYupAbmAAfXMqd0Fe1fZanRJLOxaqi
4QKl2NgtEkHGkClD7lg87P1m9Qp5Z6txtqingcfx6nCS8zmkotN1jX7z0vEhnL/19I4YE6lNDHtS
OmR01xA7fVXASWqUV245LQroBzAmgVYqDH7OuYZh58PJM9HChQEaH6uw8UXjuaoooy1sP/hfBjj6
F7rOwixKwyjYqB13u5IIVy/hAZiESVL7vmaBtT1od7J9o15nXGNS9Mg6dumtCYV2FU8hl/RSQMeQ
2vth4/+zDukg/D05OBPvS0qn0fVXU9lI6ldygMpgh3BIEl1U/4F/4m9FNxjVpswnXuT8uUOAaCRO
MptVNR0R0XvfmSG6//BQhD/0ykZbbMyNdK3VITqFK8hL59bsmMzbQyr1flEQ95b+gMJNpc2alcQK
cgxeXyv4dfB5P1asA8oKjbpLOSZKnBgbhsrps/LowRU8Aq4JYEicGsvMjPeAnVIkp6rchvJPWKW8
wYsMlYw+Ktwrfn/wZO6fIxzLyIvVEemcPfJ7s8fZJu6eYxTl7A5vG8OnSdDwy+M+4mEHLCeJ1XIW
T+AesoW2+IVri7gnu82KGNNcsPxhlQgB2+rCFNVkGfqEIAXi2uRf+OoaYaYIthJ6B14Jk0pKd04K
6hAJFzqtM8ZpMd37yqZV0HSPsPOr4HvE7b1cxa+cySfaTJaiX6HEAgAIub4aaTuPeIRyVmM8bC4n
q0spAlIXIr+K7ov2rAI/CN58MJSD3vSSAX8nsKDTOmIdO/+tsrhy+lyY/bHP7fcQRXJWkAKViY4Y
zFN8+2/OWqiBcvPYc8kzHqAxSQK6z/YQFYwMEAqTqW0F6zqqwjbLbacEBM3+wZJ3xgHfS7xjGXNe
kWt34dsYaGzU6kw731FVYkb4L7v0m9w5a4DsmfxgMj8It+yPJPvo/4MVOunx6arAEsOoXafxayfV
Guk9lUZBJRugRP9v7cWYmo8F1Oh8y+rAQ2+dACUopHGVniteQ/UzZs79kQ6qPWZeH75Ddc1aHC26
ztJJFsUJoU5AgzL4lObdZxGkhxvxmEjHib8EonQzwG8gefXoq4icYr2DLNYqxYxUqg1X73Ue0iWL
zslkesUg3MY3w1eQyJdprowHKej9xMPnWEBzpXgiNrgdBCoOagEkiOK/WE1wt9bOBhV9Xap2tHCY
tWP8K4YkD9W2uK/yUka7Xuhhb87wZv+mNxaSQD+HOFOQ0Oh60X4oE8WL0d58JJbR8O0yQdRtWqxY
+H31uqbjQJZLlq2+hE+AWTsZ/wJ06UWjB1FqQcMLMmeTT7647mT6FxTft0jT+sjs54qFEJqh+R/c
U2LyagnPtITvHyh/ujexXCgUA72Jb7T4JEUZ5VGrCTQKAi1pkxPfZppJQzM6JqtelDUWDYxgUA7P
LA4iaxQX3O1FdxzZNw3Xumzp2V1GXIkTJDng7zdnc7P4MrW4+tcS4LTxshEFFkIE2Jf1WVcFlHjo
ewVm94yNV/XI03qtMwo8ARU1yTlGI9xasnWHtmOgti7Ipj+JXJeNxYuX2Rgby9VEcv00IstY5A0l
154OQKfSOydaNbCdq2N97nYuktC24h3WCf88c07rnxO1tyff86rIBxCHtkngy0bwGrMi8qgE3//2
WFE7cLXI19v/kE8f9h/DWjm0JCOH2KF6e9aFuTXxKRb6fs6uwKhxdBcGeBoumsblLacfitTrfQbH
fdd17TI9UebSBVsHpextZVS0PsrZ+GIjWXvdxnWtahX/IH3vR0xax3bdrbxzE7eZ6+GKGzISI3nT
RKe2CEkL1b75BoRu3oVy9UD1gudbuZwEEYJaZY7UIYYWjIBnKFYz7I+DkdnssDrQSnPoifu/kFKS
xRObTepBeiqcwuxPke8y3ZH485cEa+Kw+iFKIrkaUikr29FOwNDZKvKhPg0RbMSPptraCYJb1/jt
EgbpOXht4Aq8gGaA/tgz6lKa2aql/yKDRwYBEh7NDD4Eg7JyOYbPJfxkE5af2lr/Pl+8XbKEbCtI
GWglHGALbbXQAHEKArIToixWlyZQdAMVxFQqq2giOaGccH/L/UoSvVoKY3QK+ZNtMNB4Mumxc0iN
xUpD1LF5j7x2RJqnwfNQhY0FAbd6wROCw0W/emjfPpiNJap2F8hYfwnjNwMv/DSRA8Le46FdGI8m
jCZd8nrOCDyROcUoAHwUMI7WsR8GyZ4WP0G5eswORl6yVhbbZ+1D0CWXouZtpLTRcRzMK/20EkXx
8y0Ldtaxmu+iTNrgmk3mzngkBNRJ/J8kWXVehGeC64TNUwkudgLu7p0MR/LsH6ugd3B35jOwVaD0
JwGZLXMW8arhuCkM5BPitH0mMfHVKUrllPxqpxLJb9EsrfWXb0weh5k7xxYfbqpFPUCjiQeiqSH0
A8ux3PICrCQJ3vIB1SQF4oIjs5x2DtFBAlqmq5VOG1mYQUB/M8fL02XlTN/ebp3DZdEioV/GSDSp
0w3SpkJ5v8n/TCUbOPOiG8+fCpSPVGknIznPViWC+RXyRGT1HwVXVljVMirZld1HtECSrJQ2GkP7
4jWhlh9BWX6Vf3lBhlIykMkjmPYGSN3gzsFtCKj7i6lk6fscKqr5A41nL6tmFxDY40paauO9ntlI
fmdmlP6YkVu6mDRHI5MsAE3UKLQ471wBcFs079QwColPIZDqT2Gr8mAMM461szpW2aLZROsPir9F
aJvE5IIEfEwRev6/INRx5sCEGCQd2CNjnX9AU1aeOqW3iEQgygENvWz1o5EykrQXxKKxBjqWt3Uy
ImskWaqo4PYpdOcAnQfftdUkpdmuhRElGkl77ON0DiqfBGvs4/bpxhiJqwNE0ru2uLYP/cpYQFMT
RR2nLNhUlnyfB5ottFPmzS0bDbvJ7Tst7ZZByy01714/xNIFkoVtHtWQT7XQGsSjxw5Clewy4kFJ
MLnqqyJVQ5s2lzMCZb7zZTgce1aR6UH6sluqvms4x9Isj68z5w5gut9YM0AnNqLeyf+iwk845ola
zxlYsvIXQMciwoipkvFlqI17MnoYYkAEemxfbot4zaEn8v6gTZO0FopXdYIaqCx3cb+56Gqcqcuw
gVgZt++NUJURk4Hk+j1RYdstYCsDTQ/uO5BMuCWdjiODkMXscz/Zg2L9D506BGZX0xNqZ+XNXvmI
vi18SoOaYrcdFJnbCB68ZqsjCb5qOwWfIUOEEgVPtUR1SElHjNEfl5zMB6XLrPBXbqv0p+wGSUc1
J//Bxz1VeMRxmEqLHWldPgFA9KOpasdWtsUv0pY79Bq5J9piKufztv8dORc1cy9l5QFXrah++d0s
zULWlYi3gNuSp9NrW7aoVNuuDmaFgvwvVspTz77d9qlenChxKnjY4Mi2eRJPBL0jfF50la1Q5atN
UIm5+GIwbvYshpthxuuaVWxwJUd3zJb6FrnN6w6vsQ7V2+SgqnqfrSSEVm+c+zcQPglT6VmUGrkL
hCkvtVHj645DzGphSzfYHPEC3ScuuNPceo93+X3O8axNtu2xopVPKRogwe4XNoz/ZyCI/LkoIrVA
RaaWZwI5noVw4G8u8EhLdIhcYFezP+KDjv35VKLznO8mg0uy34Kyub7hbgpPqGoL3Z64aeg7xqp9
wBaChjzXJx7TuLVpZS1KkrhZiNLsSKOSHk4vRK8t2/WbJ14e7nMU7QlR5K/TMGxuNcMZZPuaLp+0
bXVMh22CdHhOaxwa3xZ64IvNj2vuOq8F5p8gdqb0Ii8404K/zyd040SQCDWN0X//HeK4TBtD9wa0
hOnmqzlw7yyiwKTAxCXhc0HlStDcrt3iDvu7DKD9brc2yOUIPsBNYFeMPmwhYiIUQnpywkna+Q2/
XhV9/AfNNA2IIMHW4RsOhfGy/Gidu9xmSNoKVwFnEfqQSMHgRh9VrZSbmHMxQwIX+m/JFyBbS1hq
afMrQL9W2c3acPsKRohepPw3hIXymD6HlTYDifV3PLq32Gc8Yii3i8WH+3nzYibY23JB8TwyYUtx
dz69rJ/i2/4N4G3uHblNGQk/AwwF5/r7wUbp7npyAVWywqIwQng0HIvAzKe9ZZkg/pXwDVqV2Dyo
iu6AhzZ7S2zXr6mFFxxjwx6NX+HNbr/SY7H3viPgI+EAGOj+k1eRasCLurp94USpnGHkw1jTl7fp
/o8qminQsUymruxl1CtuAl3FpHxLv/2gd/hSL5QRaS4BZayEWW/Z7MjVAtXsn5h1D/YyxSDNZ3Pe
n/udNqq0jDmbQVx/CoNEBtEcoqi6NodHPa/VKpZtGMLa6lmkycigCOraF00my8ynVu6B02Z3Npn9
3hJMRcR3Xx17tIXXLuJK90vVaDQdnR1gAvFj1c9v+GI7zHR/fPh28tDLTY4WfgtdPPGBzKCWSk1X
NQ528YyesgG24ShqQxGAQ+BJus64oImxJ3F/itRZddRCgppSYx2K0KGK7Pbd+pCb33He2mUCLMK3
oCSH9WQAkMuvgE70ib/xqfgZdyx11ogl2jBVS6XEujbcyCMOPCBoY/2YcyI+2ahG2OssZQUacqRM
i1grwVnC5ZsKXeEVLZ09pdq8Zed3nPJug9VHv0zixUzVgJ2T6WBlIwoORijSKq/3pgfRIoC0Lqj6
cBPB4Rv8QJYarwTOXmgGtwKD2z7hOUctDUP7nTcJ8EkZnWU33iJCeXb9Q7Pihb7NIyr3Dyl3PWCJ
11iJcJDfzjaz7GIu29SUDIQDzP6zMo0WsL1m36xzQ2RxjmMPCMQGz0t3o8odUvfsKnx+V1ZkYFvA
oLERm4qSmFgZ2JVavjLfQtNZzKwVvHUwyVzaeH8z97Mva6EoL8kxlo8g7C/nCdeqWyXKsAIFMHi5
AMfn6vFxREifsINEgWTP8iwR+v7hFyiAEjSq1zBlBYF1ODBD1tHHjQMmrDjI4WpBP5lWqc1NblZr
M23E7S5RjVn4npzTqMrwNXbRK9jGypwQAl22MDRZBp81LUMEEa5qK4f/sucTohJefQkldXj9zzVF
iT+b5gQSkxzQIeU8n2Q35eEOQ0JITEPrBISrGSLBNWVn7zrwl6NwVvJe4dFSIm0m5CeT7CUBjzdg
MJk6ESwk/ynKWK8K9RlLzt7FMDl5+2/08EaJz6O3AVo2UcGL4PxU3Jari43j4pB/EQN0jPGpR13n
oiGLtV46j5EH7LXn8QbyBPfRjN0xO1pNDXwbG0TGguUJ+2re6SFR8JtRG2byZx30tFDMZJcDbabD
h5yGOkYoF6rOHs8dXJQlmZVIVfIjsUaPzndDvVCxt+AsyAAdzNdfwvY83AKQRsDd5KuxXfLGqqPW
hKAe9UjR+kzgu8IbvHYIZTM3xmYkngAQUdE0o2giTFghV2ocNKucWJ49ANMQ0G6seEYghUw7daNg
MOtllwfD4Koy6GIK688K+voWi9+jUSjS80BIj+6SvyC++HPXne7Df7GQtMWmeEos3ioiYqKpvBb4
Ag6MqfRk4vNHvdE7o48qf5AQXTjmThXZDr8HeKIkJfXXyRRpN2Iwtpa4wZhLDDNPyDJVuHrtne6W
X2WciZ//tRfS0PTSr7I/oRwMGe5WoaUpIR6MVk/x4wAiz/aEMiylv807qQsr8CPoc8M93xmBCidi
+4otHA3l5jVEbaww5zYwTw5mV6h2ptiQ7wZFyaE7SxbdYJbt8eugem0ivK7bAbNQok26Duyrti/Z
y9J5WMZJ6vwU4kt4z5Ecm196vhBX/13BZ5Kj9y8/dBg9ACBmwLz/rJjWR0jv3CEE4PeEF4h7/2T7
r6bUr1wL5WaQeiZ2O3sU0ckFzBcYZ35SfB7+mcC+4RX25m10u+FUy4ddfD8uvrJFpiahDP2aBOmW
+ppCpllYEvneTMBjlDgDtx/xN4H2ePXir3JnZRXFaUJTc+Cbf6z/2rakqXKH6AVigBSR7Goi8Fbd
rh5kRVfE7g5O9LaLInuhu19TzRKbEq+fGFQyE9bFQc34SUtgxwr8P5hgDLu5+xrWPBjiPCwjGUWY
bohoyyPgvdSEO27XsGu+fo2vbNALgZUmYQ6SwDEIn5sygVTiFPTOCoFkEwNic68gYnCda8GeJMJ4
TibeF1jrQAUzMjQ9/lFFToKhjQ3ddRbBk0FCF/DcXMYYcRJT7xE2+4kh0uauOjOGvoiS0XpcCxdf
kElvZdTWtEE8xrzo4hhu07I0InAhQNMqRnDljBcudD9/2TWsAb7cZPMveYgmIDrSrfVn0YBBnHSF
W4/5E65GYpzAj0PEWorkOjch/qEk4/E8LGJ2lrqsRtDkv0TppJBYch3ZBTm7qSBJLybMvYTu7Lmp
VduMLpuoWeNzY/YviUJCDMnG+qs9q63QUkjWO7+y7osQOgHgms0syIRbPvGMBqKjbby4fpUiE83A
/7BovEyBgxj+8vHyD0O715bifvTMoyWokdccwgYsUhQIzqd5LYy7Szf60RFO6Mc/9gR2j2OlWOhj
QEWokh9/1JK8lHWg5YabvkClgE7cNDNmMPn5ioxDDqaKwBzgsGeedeona1W/U1K8VdEgbYb7Asic
zqdC6neBPPtRoVLBhDh4PlY/IL+nCdKSaZUIqkrU+qqJN1B7NTvyiWXdYl8+AaUyG5QeVnJXWnqU
QwQfMbGC8DEhPuvHqCAvzOn8HEUPWDN3itOIK8fzH7a9zurXFgVYSOk7OiaxMRryaLFhFQT3HjEd
zqYDCH0Ca3A26ZButoOgFdLYiETUSXFwSN1cZvx76eyPjSfcHfJjtGeh7ryCQPAEfUGuwAOSPgf/
5DUVRrwuTqi/kIuv3yb4z6HScjUvZtswfeI2/qYmxM01sZ0RO2+HghK3noN4APbEb6YnGlOMiOVJ
XR/dx2AcZ0t1oiqzBZpkky8mxpCZ13W+IfS+eg0mFDwc0qrdOfHkP6dxxhnhMRaFkRdXBOn6N2MI
lk1FWrB427E3mx6p4d3jH83B04FCq35lQIMm8X4IBj5I0cQJJ5HZyDKdt4fgB2rpwzOdF8gWNbfa
rbSabnun3pjN3yxWLqSEpWuv7Gttw/z3ugKyWcSmDtgd+Bc1nnWUKX4JT6MH/2LUUwXPleJ2/acO
uJP9O3kPB79dm96e3KJTW4oIv39OybCxiLLbauNN4yRK81wVQNV9azhqAfp/j2Dkt4Y4lDN0gWp3
Lzaa4nXAgke2eBHcbf4kFbm7dqOIoMohfCnUn+w9JvOX6zkmqyS2gwe0oRdSZzLIJrwQmbLhdnXA
yCOdzeYMi+QAApeVf0gZuh0qIEmX16Rs0OGvU2pkmuAUWKNGxxkzDhuax7jNJuyWNWxqQrcEBLH5
pvoHtek/LEmniH7ET/wpvxrR917ojINO6rg4Oj/nH4zS5TsPFwXE+iNKM4dX6ivX2fi5xPI+znQE
d7Rqb0QxtIQcdBVWdpzNueRTyaU2dvIk+oPWlnYpueVxc5+e+BnT99uiGJR5JEct0IVMeWThj+Ck
KRmiK2MoszSH+sFhWzVkpRe3Ft1cpUAdpV1mcg3U6uKtl/RG406yTevOCilI5EVFggY6HitKzBRE
rTGw0keie4QTaKvnJMBzAYympePIVaJc+USCF4xVqOB49+dzanN8bCeGHepKLK2HpY1qNJH3kEwU
us7yhxxaG2+0SnTlLBYpbJZ8uJR1BAD3MoAWq5wK0utJFbMgLc4mJR8Tcvq17wZWnSI/Edmei/g6
20SJbLIJ5WfC6osjMY2e+LyB+UKdmgKpMrBttK4JGVtKDyHd5FHhkMGXcCysx+sBDa5Zq9aWA9rz
R3dfW9Ozhw/zMa+R6HyuBjXytBLndIbugpCZkSha6JByVvEjaNNct7vPi9rA+71D7ayZdmX/9xsK
3svoK/M3lDbMncvvHxtWCvlBT0o4BKWv9PkcZ1Yj3xIYl1npLxSB+sivDy/wmlCvVkqP6/Xp118s
z5Oexo5FDg48MwtlysMmFjGjdt0IhBBDL+u/xUum7vx04XSqtP8MtZoFFltB+/G8tXDHYbBxfrJw
hPUD2jPZq6pMywH0z6v1i6U9ASu+2vD1KtvLvq+/IfCGiTtFzinlOk3cXgBSCIY+7xeokozWg/5T
F93WFnu9NCOdBMcfvlRDPz7Rp9UWn8vUX1DR5fjE7rT0pvEXrYIIq5JBH232hEpdKlN5zl/mI52R
w5fzFpGS1pr+OSU7GFmBWa6WT33xyz+7XhqAQDEg8cOFpJDLg5UQz6FMmC9W9BHvH1J/wbst4k2n
8ZHm7fqUd2rBhiA+yGGSUYqIt8IpoR/uED4Cs3jJ+rskbstHIb9wbIaIbztIBnIieJViIy/YcgGf
GyxAjNrY02utg/YjzgYt1jvBnqZ/nBV0VmmcBVHK26dTNybyZT4nGauKrqOUQGnIQ6bjYyd3RglU
JCG1aQAbU+iRG/w18q4mBI2aVTp0lmEqUOUieO5p+VBoqBnQNFZu4ZgsGUzMYDIZGb2jYoGso8y/
2ngwmmjiMp20q9z3NkrbS+KDe9o2fkjrqwAmYWQcw+UK1xlkDVsDTi6zbhivFZHkD6aoWbyVpVkc
XvNMcwupFq5fbeyNJ7e6kUBCXjc8imQbtFK+zx/TkfruCLBCXzcTE4xcJgVTDfox4w/G8JLMVpTW
E1nSawGvnMsp14hE2VvODtS+tX1INcDeUkiHO//OnewW8rHrFancO434Dhcni+Uy3zlpQtGudEti
XNirWR0aUjGBi2iV6rsID0ehsZFakZVLekW2+EZdb3AMnNu+0ExncRH9kLtaR45KvQTEDiiAvXnB
xVQujhLW8mhwy46AcKPBUPOzrS26DvGYFZAPEF1JnFWHatPJ1jphwZvYM/la2RlG5n3fgKbka6LY
62YrCC4x6+zSLOUphXO/vTFXpokEu6625t1IBVPOSA/cBxnpH9Ew4pUM8th3undo13fSgzWFQgIw
/miOw6BWtnUInxOurkfNml2qnpRLuzxLny931UJXzmOc46CCsiKNryrfp+QAXTe7HJekLI/+kM5g
ShaHkNwVc1wRSWYuDEFRzBXcKiJtOvazW+pQ1FBCmB2mTamU+wGB/Hl0ViB+NAdt/MOBbBWQJPiY
m4SkQwNFpzWOfaPZX48uvb4UjzKlILl+wwDM2BhpYzr7qy758rlOG8bVdsGsZ39tsbXmc3OTF+cs
Lxpe/hfFuJMUFef1FluNuNNlIFtC2AX9k42wJhXl7G558JNBaIyJvc1+73lZqxGo1BzdYWQukGdA
sB2Q7SBZ5wgXMyXllH1Y7vAf7a8PeCna84XkMoutX5H+NmeBMoIvosFKB6fsqy5JCRS0dWXuo8BY
bTo1XRNwE0wbRn9g2e+sWrfIo4CvONZ80domNn2dhlnt4jatLK7lw7MYm6jKgs2L1Yy1dNj7KqR1
w569nedY4gKDEjAiRZ9VhFbUTzf8j1RTvToro0aOhD5oiruOJtIrtoalv+3hd6lXDiSQt7pt8aB2
+WCqIcK0NQTo0be+E3/eYObhu6kRIss9qT1l2j4ygCsH3XU3wTMu3mua1Oe7XOV+jq1xeTyTCGmj
ZC91rLqpMZMiuMCji0zZH+BSla6QRdDhJG0dXq+oRodplhYkTR4pF0wfcNJw5bXMIImXkS/gSv01
dcac5Jv9WnvHPLHR+lY0BX1yrVuhhlKPwqdLv4PKCZ5VXdNUXGccMeRB3Et5/wcOcyQDbZNp83aw
/2wnP4WoVn3BzU3w/unZn8NuL2maYMH42OezhWFrBunepuSCyWQ8EiFMBs//Huxopnx4Ay/6qjS/
qIZ/6/L5Gibf/teloMkCrSWZW4DA5OJIY5YxxrW6w+po7aN6Dczwqg+WUpwrqGehKQNIRJgMTxgD
KhKI/y0337FkPMybQfSva1nHo0gSu7hnAb5Tlpzai6DZfOjZklZqSj+HMIHFYvfIiWoyqNd7GKYd
CMweixD9V+zz9rcxnH4gLR3oilo2OkQXIBFwy8Qbejss+i4AC9JvLFdneYqKvqseZdelCB799907
Tccj3l1HFQSmAj15CQCuWaK93teWkq/aW+dH9KzL4Iw05jLLOq+BmBfCFHX45vTp86b3bDxPJ+Rr
qnBaU1wWPKcBt2bzTeLSlNT/WtegUnzi5D7bD83Cz+/Qoj0FPUxspdLKJnpylh8hwU5YuXkh1sAp
m7Y4y3aFEKi8OVktiMoXLRNXWnJbx69HqcgUcvWov3dHKp6sikcQROLTk4EFtajM3R3f6MteKDJz
y0T5zWwU449tpywuj72s5YHxxBa+WIHHOMg92Wh/HEOy68v8LuvZ9TgobhcVSXRo7zWSZ3x+2m7r
b0TtA9Hk3JtW/J58Wl2nbWX7jQcmO6KlwTw2iw6UN67bnnaa5LAwyJbeh+EI1zqw+IvWn5f7KghE
Z9F/rKXdtdVuk4a20n8BD1TsifkL2iy8twZDfZpOzbdbmbAeglwaEZGW7e4q0Ht2O6v+NPY699xt
7r1TIIUbifqYP3u7FXxU47w3Oxp1BiWQadRfkx3gypnV8tokRrzBfevb+qwn53S6lMsvKxJ2w+7Z
Dgimq4k/+gQdQDLXfN60aztSw8yeCjZKzOG8UHaEp4djK/Zul+2CSKaOHgbSGPH2CcuNEGukbmG2
5QRuJeCCxfgIJVI/x2wzXwWx4U3iCSrCYsWshXc6AM4GCHVv05oQz9q19WoC2BK25jb5YY1/jdWd
z+1eCRL8cKbEkJrn/lK5hYReyG6VvDbsXCqiK8yfa2UvjYfm1SIM0khdFgraUXiQ6HmaDTyx/pji
G6SsEkM0VP0ZDcoJzeqljRV/YcKJnxrY67cI/pJkG4qgyytRNR1OsPDEXcPYXLJajol3YJtyFzPB
YQ8VTXl1EuMtbgo5fxaB5Oumg956kHtPIHhe+ysRvv7JV3gNSgv69baRH4DhxrcmyVQLI5f6FYbH
9gL6mFVrGdmEp4xUd+GPhVnDeJnVJ+UwDo3//vCy067VjEBplExJyyRxEvcQ80TDCxIR8xHRcMgs
Vqe9zbfOir6UvreFwugg25Das3PZyfRfLXm2QSJ4HyeovqCMkWVkHFubo1fzwDKQKCFRxAza5z5k
mKyBECHPPxHhBXvgkXkgiDTKoLGYN1k7uprePSxxkmBlIFPo7sH/UZBaQB41WuRFiLLamciLpOIQ
po14zMv90rb1yR8yFVvFoghWnpym2GJYPhW0QbBYddIwC/wbrgCQIk2cwBEXS6iGo3xxyBFfvZpD
uZ+xGx0GS4TdhJ5gVcKd2wv75WzR4qh8F3NQ9TGgGKT8zczurNu58NxhAR3IUL70qWl7XCdT2Uhe
tSO8mXzgsLNSDJGabqALIA6HyHl7q+l78YvmAtw33/iyDMzjmQUYW1MoT1vRWVrjmFunBgui5O6s
v490l+irfZoYdlU8Jf8l4hXqDcz+VI0GUG1bNAGYQe8Se/LJLKlxpZEVQ0BhMq4A2safAfaB6nPR
l/sKone0a7lmhAccQoZmrrAJAdo8Q4Jodw0Ij0UwAScftRBDpLiAptDRcBBzOv8wmzVPKZrjE7qW
gYeM1H/MgSaz9qrhDmtm0QbFT13E99mGKW9TGws3azydPFJ215wfxYMVtq6rwFmNGGUAIys4AUn1
qFR3UXQhARIajtz/Y1RPjlhvYFYEvvVQ42WYhDWAtNRJNpaZ3PC7PQuVqr6oJEsrsTQL4ExVn1W2
bkCLjHk/9Rg2umkRnpCCe/a/DIx6oW7fcV+u2Pgc/bOmJ6rtor8Xjhwc2WfcA/cLwK73jOhOeyQ4
q1h9qGllLMTF03RBfYWteBxDk3U/AQcOY95Jp4axfIkCMjHnkFHKD8ZBJ4smh+cpfq6z/1uJpwFM
amq+rubp80OkNoo9TTyZ7x3N2hTMZkSx3mtjgNwrKQRwhN7try64Ti+7QrZ1h/sDFZVHx02S5QMA
PkkW1W938rd4FfoeRXEkywsa+4LoCxVJj+fBazJOVujHuv+s2ANI+rx4GN92aOyDG2xnXFLfOoBS
7LEN7EGoqCX++fNXrM7GsSFqOieAy4xaSdH/RoishjEq6XguRXIiCPyMBLjMoPMDtFGVjS7dqvE3
e8MzO8E4Sqta4VsRfCCz9qqm4UofnfvC5loaLohX8KIUpRGVDglQwMrvr7p+AHLVevmRpahdvgMH
tCTb9ZQ5+KQFvElM45v3N9bUgKaChPbG3pJmGbe7VAzkx1dmbO5uoswYljZgsRVrABl6V6BFu3WZ
O+DASs11PPwPeECWd26ddk+ehNw1D94sDp4SiwF7QFzhTTOfiuIS/eKjb54LQtBYQz5amg5JcauR
u7PDtAT5L1/91CduuabWUAHuCMRNCS2f0/uoEntnwrE630Y9WiPoQf+Ub4TZqC47JFuwHizKwNDl
UQdNQcFQwYKnD0aqrY7qQDuS6ie6erZP3dgk98GVHxDC5Fjjg5u3KT/R3tMfAdWproXocL/FJAjE
J1sRPeY3wnhKhRr6TcBosi1uFjLdPk/s3YXWvebBJluydIXL16uMzRCC3m4nzd7Wmoq7ASyY1DUd
ytgiictw6uciD0p5wyWzzaHxr1LpYCR+ycwKHKXaR93dPViIdO1N+RBytJwsSXuJ7E9APhfIRUlu
pRHjKPIaDMFhzrGiBntlS3JtDnOqtROFLSQ0tX/BAt8rC0BUVcK+bjcuzBbZgnakCJtg0yauUxHw
Tz2Hd97/sWNVxeUwD7+OdI1WZQLRNpA6NxpE+/hK1XPOtRNwbu/arH8aQY2qUAlplj1TalpiaNXl
P7CjySfgRP5qy55G6sh23LlBTUNd8JZ9wfov/AFBeCm6rb6YvKglKqnr0d1jSJhj4nNCvVkmzYWj
YXuSlfqg7o6Ypdfvm1qz2FZMrtne6vSbUBs6TWGgyPrkA7sdHVo3fXkeVI+aLEMEdpcb0gXU/k2r
AUp46x/YXhH67sHV1FU/7dt3b0ap8fyP7MTvgoUZu/muZUryifwAYMh08PiZkblb69KkvKeXfkbZ
0tikgk5w7BUV1Pa0V8GxG4decG5MxB7D8798c51h3MpcQrkjfIRD91Uxdx5gtATqW5cdz55ynkxz
XRtTD3YpoWUh0BEfcj7KEnPI6zlmC6R1mcairF6v99IxkXA5HqnOKK6r8Ig8DsF4I0+6fx6pUPfK
riBdnoq+TdcVk0jgDlvK3Y9CdFR4x3EkShQMosEqt5KaNhdErkUMGPG1yvfun0bePYmd0XIenD+Q
mP+R9aAaiXhgY75PWmmKOaFZjr3jKMov363W+o+0FjFjcWAMheHviobzwbshD4xG+ZjumThb3Lzl
lLOGt4AHQhgY0uYN+zAJAU8Q74GsZuG01azT0KQVEMt7ajeH91uh4aISxmhPEb0CBnVh/DSiJYs6
fTRS+xpIN5/vXiEYkoKTwuzRxxJL9OfKXgm9V+yLYybTYQ6svFkY6Hrecv7nKOFs6nJpOyS5/Z19
BNKtAS5JzGDw9g1l6d5GC2Utj935Uls48W2k+L57rcRLU/DJReMwkH4uayuR5CKYgXvU48Yin1qz
2NfJxiRATd3NdAD9Tpz54vGit3LAD01n4r/3VxRQkzIR4254H2cjlY4q374vyN1Nf+FZSZ90TsyV
vVzbnwwnTw6cwzezMDpYng4guKwOaI4L3/YpT3tqSIH1jil2S+FPAd83UaF+0UcAUjwPFgUPAysw
kT3K+80geL5FLzspSW8yQHMOpKX/srEHkna3rQxmKLgV/BDDYH9rNTUgx5S2PyWbpMw7xxxi4MR+
tisw+kIFVGDnj8FeAOMrO/PR9CSfQW/8fPJMTszDimpBbn2ki/f/lOzyiLPM4kbNCOEyXZjLE/Wz
0t+FypUKV27VfzbNsQNFJhwIaQFQVoy48JUbZB0NrEa/PC4Opa7WZ1L6Xtj7aomPAgNFIYes4NHS
4PgjNurrRujLRpIRkV7OAMmOaYkdcPxINq/D//QxY/di3vATk8Wyn4MPtWTrj2mN7EEdnS3Gk1hn
SpR2Yy+ySr1LfGvx97gOnv42RYfntvmmiC+79syyH1y6P1c3JCdcFq86dcSmHI26hvsPGgfIyZ0M
Yk5N5gWtwwfjafqtZ2+7ozm+yHDm6ck1s7f5lP1bbhqIhJYlys6SGHlJqnkxXftn9ukXIGzM2XrT
gGBGfu2a2l5KZoCCoE5IdRpICF6P/2ry5PFMbd7S5lEd5bwl9V7hj2sjkX9rkCvBFfQqkFwCPm8k
6QGiw0BM0w4G9U5XPJbwA6hqp03a0nd/f0d6u6se/0xYD9ocGq0jlwV1O36M17mNNvLjpQrONoye
z6Jz4qEu0TRjZwn6rt4hMxi4y9rpwiiix/1P7Unr5w+WyELGBbTLC5aopNewIATcetMsyBkDHHvM
8VSlnzZsDp8IjGglVaDd6eb4s08FXTNIoPKov9/oTcpIY0CNvO8qCvQDJ0lRqFJR4ibbi79Y2RON
gVinIvoXQl8ANzfKgP4pJRm5dWi9tOSXA2Q7QvBJU9kprut1M9jtIdMxF3aEmjc1Ce25WWnVvyTJ
cSJNLdrqgWsdJiaIC4MfuyEbI85edYtPs8BxphrxvplBJbxZ5bioWlK54vFqE179fc3Tj3ADfHry
yIXrsdT0IK+RJFKVle5Dia8vCoEtY0J3BnC+mPYj2NOuPWmdXbSw5QItiM22ofkIx6l4fc0iXLf0
4AMKnad7yHMHLtaq11XVQqv5hKwwgo2EFjZKrbraEuAIc13ah4FRUCW09xbaRwIZZpDRNm0RIU+9
K/1a4UfFjx7HwMiFajc3C09pM3feiFyl9At9b9qYtcNd45HiTqPhqnu2imLckGoGCy3o1wzJjOC8
NZNiOjHjhICsHegmw6eGzEnkEJxwq1kS0ijpvkBPub8as5IJuH0gC7FWYp1L7oUGDShlMuI0TIlm
t1r2pyZ9mDqN8fZb66Z1gOwrvdgdG+5auORv/X9t1wM5GNrq9yBlf7Cm+DlD9J4a6YSX9EnWlRn/
u2xEV1Kvs2RWna8HMuDzPkODcsJjT1VGrTSH1sgJXSvONsXBliAUUqW0VpQops7/tw4Dl8DmkLhC
Ov6g/t3fDgcq2SPACiMT1X4zu485lIJLQd4uwFY9VyiggbsoB5SfZTk/U+llCFIQesFv0vMv33kI
F8J9l9zUp5LwVlRgXkSKXDQ4Dhshr0WSgoGMTmRFwxRsj7rI9oaAT2Dj66je2xHa3g6oAsndXlLI
dtm9ZzKpdXoArraBZdmRPXZw4iTETvQadj2jdCPn/zXUbIGVCQ/6PedKz62ebKmUVd7f1mn39E6z
BlpcMsZ0qe1lkMOiFU0CKiZne3nqpXT26fLSo9QlNH8hmNFlfNsFV3TkrbALC4BQVsKEfKqwy7MO
pqzTXtS/1MZada+0rs0eiHYjBKNAoqWbLRO9dTzMpUFCznn5TJ3MYyQRrSPaKbQ0bCBX/pC64xJ0
gurZfJQDoHj//Z6xj7F+8I7aXOXFkQFUn1Cz8umc6n4IhuDwmGSGdnmHl6Gu12u8lqN5B3cejzWH
/7EkXNDjbhl5FuybemKB/jFFf5pqRJh2k+4IPUEyhfxaLz0WOlj1A3wM5sTnCO/oFXxd0tkuu5w1
tjof0zaJq5HpBh/8U46nr7v0HuNRnIoQKWmCPqCJbj0buHOuf289G7vgCc9xMxDTH80B37O8iZ2g
3XTXTDziY/UDU68+qCga/qL1b51lK/cteqVG+VzsCSWVol95M8VjgdPVwa6REwEG5M+fzI2EwNz8
Qddgtg9MiwoZpXeo85Tz2gbsQq4vDe+OaBZGJ1efkjVGe4281gTOpzEWNyLNNQmoFzclyGzTeAC2
VfbhzERZv5ayOrIWPwZQT8pGAL71RIzekZoXxBQ14/OfFP+GxGFNMVn47j4/KQTJgjHc+6XUA1rx
VggwsxSx3z315UKe+u7Pt9IRBsoNPof+ts/LHUePKxMJKA8c/tFDjNKabUkt+O9a7BGsXrJdDhDD
4dCDR4KYbZCD+wrLghlGIziWj2fAZddbqpUccAMpXTQvZlqS+p8dz0zPZzjDmI5nS/gphf++px6k
pZmhc/iMNB6XAjPe0tdUM3+QdbKxqhjlOTDSOkqA4B4Fo/yTUnthQ/wOdDXRq8bvG14MSHHl7Uc+
CbWwZ4HXIsbqOMqS028bXqlFwkTqrXYaDiejpuPrTH1PL7rchOsiwgSqeWvUFgVJsuwDcjul5KxH
MxC1exEy0BtbgFVnHQPOtZSwuCRa9Ikf16mdag61sx1aPJzP9pKRzo333CGjnZN4t7TwLWCRfpDR
utqwGWpXkJbP3ryssX3GOg7K4P24LY4UMHvX3MwiPFz9q6XKU5T446Zqk73+9gBd6OnkeAo4S2Lm
8Uy2nGaHNGytROOA6mHw6ATD45KdjtZgdt5tKM74uGfL9TN7dv0Q/dDEHAT5YMOQrWhnC7xNvV3v
/djubGbJRzDp/IulobicCIAa+feOOdJVKhuTdryaN4eckOjBlcY2vp97xkLjTqfJXlri2Ne5lr+K
mn3ng0M2v5tcA80rqQgmfoMwQiA7r4Gqwojxln832AokVX6iaxXMijYZWqz+ZYyETSFvuBIuPxHx
Eyi88aV7uoo2c6zHAWS3ye8w0oIovE35LB5yFVUnNqqZAnArxXWMLccqi1OfiCfi2OOB8c7mwueo
FoxeT0vNyBkRSFLLwK8jBPILUm0u8050KEDWQYf2D/UwYRqToF5T0cd7XPPJb/NCsC8YSfx0oCX9
75ddYgusvKxsUU/Y2pu6uet2P7tEKg8PfhJza+4vrt21Q9oWrKlHvElOt4sbZf/1tkgErxYW2O4F
Ayt/MkhkV6nBS4hTOO7b9v82USQEi1Jnx8ycrwRv/to6K1RsMerDox2LfD5VlX59NvydorPKCii7
KHTf2l72qGTPPtr/XTOK/aWDHNcrJwXEd5S4ILUNi2nJRokXap2HMwWmLUNRblKRUO3cdySNT7Am
jR0iDEkghrbATPRQor6Nc+o25dPqq3V5LtbXINb+4ccnEOLjeI8lD9FzUh2L06l1OjnjmyxMM9uA
xCPTdVvRuareS6xZgbaPsH8wEWRPvb3Txc2SQpOrNtgc1XrYu20Pp/wSFD2Xk3XUYdgFa3UfB+pX
oIZewCB9MpXD4zx4RBz1v454k1N95zOu+j+o7uZR8ac+BF6GgbdxFuhuvfG4x7496Fl3wbcHqFuc
/63vPHCkq/bPNHvsBEdTEDhn4eqMVrIbVxQSZzFHA6jEIHQM4EO032w2rjrrcqg8b9XssefDkvlr
l8gJXy1S404J5iJdMpO+ki6MSFDGo7KeTUU3A09tTHZ1rYG9ydmaglFVD3DQUAGpb6LY0By+sNwq
yezBYmx4vrLY1YxVxA2Qv8p6DT6SZ+ZDCVfard6aorTeBtzjEe0L+lTJk/UrgXVXuRgCALcCD2ir
FYa6VlR/tDOQttAV0QGTE3wfQ3YjZ6Uxr+FPTJW5kMiMpkl4MDHbEZROw6gim34JhNU1Fccvnec6
/j0BN2G0NBN/SMu9ffKoEznoaQhpSjHGCsDfcHd+5WX7tLkZFLoRvWkoT+xBdm2EIAFoJ6+TfvPK
G/Hp22jrp9FsHcp4bjXAsKkJmfrF7m9Yo5cT9EgQslzJWH3WGdcq+I66AHN15UhrSdXDiyPXMYL8
N0hqVF7V+7XZM1DJd8MI7dE8BGAHAt7H/QJAGK8CdyBvvJu1xnUzRYCfObWvLUX55LW6g0rxVtBP
AiPzb7n6vUMXzhfhw1pM/A3brJm5rbZSd2S0zjFP16yQ3MhcC4elns6laCffJ1Grve0t4CeoL8kb
8wADQr17tBsCHOtgpy5+OjWReZgd+MykZtxLtSXDYgpYvoqWuTGT9oQuhuGokvLeLRpgQRKavBuC
/nu4M9lR8VBqMx4J5qFR7O0cVoQIYNN2oP/i0eIvVpZ8bhJVR4SrILS3R/WZTAxMCrm+vff4Y2Sj
jyY3X4mehypAPFg1Q4f2hvET0ejwuXA7cv6xDjgZbyRXM6wmvxx6uFgFqlVtOWTolAYWKKqFmLOu
w9/8Cdnke/YOe8AQu0dHy5S7/d0Ba3HhWlTfv+o79E+7OpmnQFcIhkmBeFfNedvQWSzFojAlf1eU
UgLAFddjLPB7KHgHQJTj0313B0xmrPMxZW0DOU93bC2uUUlOS6HxvSwfE/9zYg3mUbAoEdpwOMAX
guoSvicp8uZ59radXT/IW4anSlsFgEqpm/rgQuyMuxGhs9qF+N4hgc2mABI3mGvIeIeSfsc0Nyji
UZ9Gst0Ssu/h5JC9cB5dDmQuYiC0geI+OtYG/bIfzpnz7qKkIPw0JluJncODqzCNcPryK18jREcZ
MXBZeXfn9Y6wcAnmXxKSnY8baHWgNIwnCEWJxcdXsHQxSCpk6DBtQbe1PvxGtFhPODVd8eBG/+R0
akngVrm9fSjqUESwC/umziOQzCqSElxWQza2IhysWA/s2kmNleHKPvqo1e6sK+GKtoRixZafCu4A
KAkv/mBct7eEjda/uI9iX7R8J7wcFgnv1t5I57H17I8Yc+EJTMTpAUuNziGmQwzEEaoJJCSSupQ2
r2i5QD/p768ok2VReyWGwGrMwkqCDsKyGGPAx4BM/UjHKqf4Aqs9NOAUK4bQQ6FSCKDLE6CWDjj5
ASnK0hOazIXmJuYFLZKxcwvUFX+aZPW//z6/9ksnDcK+4uY4quiq2dKC8xmXCyWYf3JmFD3gfcYS
5mCT5iw1DALuhBSTitFsy0ZDVVIYsmrirtt3bG0eFuqxBMUcLu+9i11TrwHlwP0F1guUNLi9tyer
r7zRWTXfuJTBq1US15YAEbY5HYJH7lk6bs/n08o/JjYRmMJO0z+GGnRFTqFouRFJnXj1zxU2NNIo
NGDXwYKYwLG5L/o2XOMln85DwnjmNXUl0UxbZb2+EwgsXTEgBrOfjxr21toyHqfLZgT5VLouaz+a
qQtcV7g5DBm8Ffr0R/CGS1xi+le8xrSKKo/+FFBMbF7ux1gUeaomvezpJB7wik+hoGcz6vzE2FtQ
3/ab71R+O9q3TDKnRcSWhPo/jMSUCXtt0kFMFcUQInKV1bK4r7iuDnt6Q6nYnjcSb3yoFv/Z8JnJ
zu9G/B6L2HrwRPStJJTCRnQX9xUMeQ6p5mcd72VBANyX/FWyktbvvY4rBWjQUYF3Osbl60DkcOEA
aTF1Ylu+/bhRJMo8cSZ+QxWdyCDDb99c5ibIVhhGZHO2VY1OVlykFO78BaLfqGe4BpT7+/smtr8F
rFcpfNAaDDRC5aJbG5mFgajvL4noD1ve9J45c1qPgBp7JoO5Yojo2ak56LOxYHBnrMucbe6OQDmt
QqCnxWnymRjmb0VQ/mug5JvKNR0V/BxmzygGNtg3IyBR23Kx3GPtM9c4dibiqPJjltVxh8jgbmri
AlTAb9Jdxo/46J0I2eV0B4hW/IpXiwLV19mv1u9c5y3hQxcsZ7pjXMiUqSZ7uMnLZfDYyHlEqmw/
UroUvT3nFssIqejCakaIqTmkGa5AslHdy/0/Z3Cwzf0gsnCIjiPiRESxkN9OgFgBijnL/iYpbJR7
EU5PP6aIiT4Rze+sswDjFh0vml6wToXlAsdaa2HkED1yiFBGvkBFYQhV4WbjvDXXaXtCnupPcYTZ
jZEQpW5YaHev5lhzHfWYNbAIUzLfRAsc7Top2ug/ncUajUfRuKKpho9qhMGPDi+shzohDo2NccXw
oVrJQJfVCRyJcOmQvf8YfiZMmKEtllgmT52Bikgp2sCpAe9ydnVGqxfs2moG/BC4rvUiv1HLfFPw
5GHdPUrpF7jFR1DvJb+JzqMJ2tvRVuFNjNFZHbVXWsFGlZTOW5JBgAFmUFAgLPM7cKOPnLtXXDad
cdKbIcJfGD8djdTRYI1oZKK4OjYsrz1zZuGGCc+SsjKzASxxioZBSA6QQPucUU+tL1x/W91eeiSH
GzJIH9poOW6v/1qIHvL2REGdLvfxS3qq5gpbwr9+7PPiCZJ11FBojqpyqpLAvfK0P8MuiiL0kuVi
erNjICm3Pfir0WhGF+4UCxsmCNputIhcjTB5Yc0m7zXMKvp6YIy+aND8fFH6NqP3iV5SfbAhqD8s
MEyyBodTuBklEG/khwQrIQAF8NHgtcTJrferotIrR7XND5ncfmcGyW00Ku2rZBaoFAVM2oRwOtnq
mHUPWrrGR9eQgGZXk/Qw0QNlWjNPGruOCRegfDpThx3G0lZu3LJDepNZjx99PmI4JnfybH4ZbjYA
MW+Qh0GaHvnNrptyG0o7IOlDa4/ukrDPCs1CzcvZjGBIQh6Zc+v69hAL5tM4lCaJBq0Y8H3OTgmW
28q1Nv01IDZ45RVX5sqk4ahDNAxOChR0c3mjNHxkXBXqSqbSWeCCQBLpDa+/riW2ZsZy2HYRU13A
7/JF1kB5i3Qut70+W0RRDDSK/H2WAvEAEXB5agWIxZZm2A/AWMLTBzmyMpcrZye1gVDDwQAEF8+q
uBXBKSYnpBrzB3Caz3L6GmItAL27D9kz2HqOqu2Le6RQKQkozs1HHLc6PrZvh5+KVMPgqXXD8Uix
2tfE8ll48NSs8cqoNELtC+ZhG2MYENHqxblK2q69IriafYYjNWD2tKlaQWdeC4QJw6J/leH/yW28
VHwBo+QkPKXQHHIiuY3v1MhtKa8uYl+zna+4yxF804A5/dEp+q0qPlhvRIV1SRCktEhlpmO7NDgg
ArwgSZVjspSUCQaa4ooXqTZiWV5X8Ie9MGbaTpQWAGoXHNYyOGuhYDhzSkguHwJF6JPNI7P1LS2J
NvXaJbGeF2t+iVtYcNYUH2dqD1ea0yVkJyhJHHfBlloTHSWaspsaQ9P0FNUeK38IPtGNAVDn4Qdp
BanAoUkTpr+OzTeAXVBb8mfAP06FbeEfX2sONe7nGSYl/uo1MjoPgZTgM6UXrtBwrcY3KUaRRpmw
ectM41uRuz/QHEH95+QCkpLYXwBi8SqUoemOxY20eX+41FoSTtYi4o3qNeowJyqAVFrgWlZreVfQ
P1R82GbnfLHb2UXGbcIKfUIUqZ1vYv3C0bjxjPzwt2nFKVp2LOrbtDGlaNpls1/Vvn4KxZ6hghVH
HOjPcATyJEgQfc46IZANRYK26z499HR2zkrXA+78zG3EegDJG8/2ttBSoXBjCFU6nHQ9dsbMjnqO
HH9ZVQYap9mqrysbcLOICrNT/f5dAtZ1mkZk1ne8eJvYS7bcfoJY+0Mj08XWf2rKfmuDygU+OKmQ
N+PGV1ejZLMiBJQftgl8FuGuy+F2XapWNoo0A0Z7F8yUnb1E1iH0F4HREjkqXBptp60oP/15inRX
k8jJ1TJJU0h7VhtW6TY3tSv5wdKJ4eu8SDSUrBDx3tplPrbhhvB40aJYMFpXrLFYv/5FJjLHFB8R
x7tLZtWYwWWp4NGPd39xO9WagoS/s93CaKnEI2czV3l7+JA0vQb7CsC2CHiDLYpX4TpJhWOqfm5+
par599O0358BNYT1u2tp1reS/ktHnS4Uv9nyjbz0ncd6PwIx1vNNLV1xmTQNNdwLkIh09wG7QWhE
7H0hyq5DNGZTpHpvuvh/LmKUoht23NZNsdjQ3ubexkiBeN/UphRDpVHoa6xcpk53VS90r7NEhNKF
P3InnjNTsL8kLUM40GGiGgjTcWkljnvMhsBJ4QNrkGCWRI5GQPf2hHIa0bEf9Rz0mPdFXOUWr17L
z/YS4s+m9EFaHF7MqtCXu4VVWbOgxvEWgC91jGxzQnKWDOMqAymdpZ3jxQLE0F8SPWzAVirI8JKN
CRRD6KMyQu4jsKBOmrWPMBcKRF+sJgJMeeLlxxLI5euAw++MdS7QlDvdQdYzrfQsLUMqIdI5lcHK
DqYw1TxOcPtEXxpO0zv7Qw6qUXST3tMkxedGZu6DFYVuOPkjSgdTx/IugmKwoBOugQzx2TRDmecl
KwcucbbEMb0cdTw0C3AnECTliXrRgzuuYB7jKwT0ghEn3hn6KXLiF6gK5wJNyfWmqdl94jV2v0wg
s2GKj4Oou07D6XfKRdr055afx2jB9jEnMLWnzF9pB/KJ9gK6RO8bjLzBzrMbaVZqoZq67qhtbGZJ
UPMRMmNNGJPH2RUulRR4AuXy3BMRFk6IeJyCFP37gLcOGBswlmyOgiGsJdXD7s9mGalaWtuRsn8S
2/q/xfxJ/D2fE7IGMQ3n12jEsbTV2KuTEB+W4oCobgPo7SZfv9I9QM0KOty/0OW4484UykMfDpUX
iYMHiPErpZskdkytttxLZRtJhJoCi1Fx9RXeE1XrgDQ58BMZdh+48TRhkNAEQc6LJMx3LFpowBa1
2aO51MW5fKrp8J4jK85cSObNDMTfdF1RX7zJqrb+r+GktLdaoOujXy/HJocPI+FL4FIpMQfvtbBy
kk8yXax7/d1hkDcMVJbVdjf6jPjC2BHOMR96z8L4CcR2VHs7kLc4xmNJa42iBR5xncRk3hqLfaDy
vrOUubrAiYjvvwCLkdcjRFmCxcW+NPL/dNsbW2hyOoviBerEnE4fBhXRTQdddvHgXc4P8Z4jqpPS
rEKkKS4H1TB19jOOUz3Q0kYFgl266GCfGentb71W2SqfIcdiiY73loQ0/HzvQqE6tpGSsMUC+Bxv
VGvGYVs+Z+FYjOv6hWTQg9Wv+LPuSSWUeHit5NmJAZiXa8zQy9h+hwyBUhx/Y530SBWs/xpZ3Bl8
xxYIRhzJbyLfnfdqUY1oBIhjAsKRF51MGy8V5p75vasZM0qLy9GwkTvgP1bc1HuYA3NBYxjsL7M3
k6uUiCj/oX//EtatTiM6PfwBv2rRShZyUY1UEgWW7X37Qlutfl+llrfEPe1MVyB2KXiZjX5spB/K
joGjg4G6JYmYoiRuVEFcVDUvcc21JMZIXozFAvrtFdd4I2L7GUqnlxUkQAQ+FnT3jbBdOZALHnNS
u25UtM7jd+BsJf1ytEP0qSVMtHAsm/ssXdN4D4AQIqTRdG7yDSEl7AMbklWux2spErw3s3d2Y80z
qM1SkHNh7AAjIibq5j1G19cT2gpo8BLDtFeyYbjdfVtZRPl6jWw85rG1+PN9zQ7Mk2G6sCgTNZxz
eS8vyBwlnJb76+H2MikZrfN5wg6d0/YazRdLJTcTJKb34IxWfWE51Tw3awsnjDuxowbdj5SQBvZk
tbJIVw8PXpjcaTTONdbF4beQAYEZAHFjBeFILZcZhc7UJAKEbWEaGVlKtoVDnRlN6vm9D02nvqBN
Vd9MA+v6MTCr0gvSlUzbswNGYsIGhnBxVtExDjDx2qNflfxbOBovYQBbCXIzRgzkq9CKLLRyucWI
B2BXKg93oYSHPqrsZ+vUcQOWmQHKo13YsVrg2cVyxiZytwQkkPf2seAmGZ2te2htutuoSITcNrBh
zW8yQTGfIaKOevmBD3GWbD2C9N1WWBRGIUVqshOnGnOQcOUcjTb8VvmJscUvHNTv7mzwD741u1Ob
sm/pIHEr5dW9292IcsLabokogGUIGHpHzu4Z8aYd1KysFUKHB33iIyX05Hp+eqhbBP0R045Q06OH
0xTtxRMpM6m7wAv0if7lbu950+lXZDqPkwOcuVVw7azTcbHnkwHY7z0QHa8GelPKmhXne9q9RkdI
P/PuTaJ5ZQhNcH5IDUIT+ERgsQOQAF1UxirKCWc2r3+tIFrsv3wXW9txc7QUFHUHcUd5kq0CDJSw
fdV24yyFKdKaWdehWt1pTRZOdMKrDfdeU4bT3x88SE0GnGsrAERnvy1THtfB0zWejInkR9tmLTYK
Tw1xIcjiuujBroc4sUKiOmRul9+XDLzYv/3S5UCLP3QXRizSJsHeBPKPqSdrIVlxMwu82p8nNADI
7tf8IYY4oxouArJ9GeX+noZ9+j+nD7nfLJTt1qwwfkEAsPbZyrqjQbvExYImsUh4EPbOIsPmOwWR
Ej7H/ZW3/eB2WWIESF7XCS4xV8wukmL68/X/lv/mq3Xx1opOCQ/8YmrXIlXmhsa1G1yFET3AjwkO
FZ1AXwVW4KV6dcE1GYE4F9TeUvMVcoZw54pQwhNKtHprU3WzpSKlwfYjA4M38itdb36IAJKYzGAp
LLtOoTj+MTKgPtX83fntrqOys5HP1v62GvoQi1EbirWx2/5bEf+t3BgMrlX2Qor9APDBGaDLsAOe
EQbvbvFtM4Lqcv3vSIrGI/s+/+LBFBIwFjNwWHrDae6r5iTWpfMx2+9/VSb8pzsYy5/gC60qEIdH
JMj1HOJhDGYlMRoWT1KbuEbfuxsnQP2uBhT8FhuE0/mhTGZRVozRbjVQSCvcEU4Q0OQRSSw1M8ws
pvZTf9D5lJcpQv50/B438lJk1MOOgcOArF49t5NmHCw+7J9wtXGiCUyzY5G5CLzs5kS/9w01rGoZ
KCCDrhHXqLs/y97jOe19We53m3fbr8PcaL8uNjyNJkzkB72iYljkmDR7x2tUbEyZATKVlUgUvMhH
Ji+99vKDliv8cGj8jY4HeqOWdXTXB68y9yD0L6x2h8jU7MEAdiSEe+YssXI6ibywPF2e4Ky/aY86
FhurRMs9kqfkE8sj1vOIRtwQJ0z+HHC2V5iFn0eLL7LVRmxJC8psZMBsC6aGMa/eQMpymgGEU1OB
BkuButSUENVI55jDWKZXaSNWysSW7tnGkOR62Knq4Y+HBLCrcStENVJR1CBmuqjdYnVtJjPXYARG
SHcXinp9SWR4VBgDeEWkD2XAX0XcModyWIrZlJt9eGAfvb83Svx8+LRPUAoXKdDKtLbsHb12ED80
rz4OIVR+ez7bn3UudhvBBgkfXZzEAGHZD185cFln+hTAPCJ5msRPkiaOQV/Nyz9ZBwGqOW0qEtt+
ztNsLpyBhBVnUdwa7qofQTBpMGWldA6bu7eb6tWVLOn+JYxafJu1VC7xRtjKVoqdNd5LaDdinmuD
+BVSvbTEgJKsxJvhGx6vdQGLe9RBT5GhEhgpmLVtEM3Dq9ZiTaI9JnnucYg3h/QXWxYKFN48vRLF
ivWJTirgxFPLmlPtq1dgKe+88UMz2Gbd4EfmMFCgm9aT4BV2gOf7REyfoab86R3e7wVQP1w+OsWn
ocbNAJIsHvV2jvUt/gvmgLP5ZGdLOi8Va5vuwucbmiAma7YPt729f6GxjqZaJ6a/UV3ZUCatDEKU
ZHHSaGvRh6Le1VQvWXNnUkA7hink8htR73/fNamCfxkBXcR4ge4Cz16iPlR4hBHhAmfT2Ku3cwtS
Bx/q0/Za3L5tbHykA2c9uFZ5PSyf71/y/PGMfOcckp/25d9llac5tDN9dY5zLG6VNT9J2fw/+Z8N
7UCvHaPed+naslZ1ISx+SunaBw5nSH77OCb59Zlb/cLpQBzZ561XeJDzfhjDX/qepa4uLOFwzV1g
U3r87sgUW5JMNnHZLTNX0n05E3aJOkCWqHVcl1e6ZWSIyKyBrnP5Epkm0ZixLLxW8j2NZPmqjLvH
rnmptIOo8MxNJyyehRV8JxPeIPUI5lr1R6KiO1KB4R5kFNhtYNWDmvjb7XoJzFezFkvFOWVdI96z
h3ZHDEZWm2hq2arFoHF7FDitCv09c1n7khmrZlTT7BEa4jxn9yj0aCx+0sRFrqhoK0QM2BBVFgnf
nq40WnxFh9Y+RRkoxDvHg+UQs+tqCiuIgbJPfBhJaxbI5nA/Nv/5kWaH1mb4PV+c+85AK5z0lkrt
noKSwox5e86FuYCzdBfI9knNPURBqVc2cmaauFzAh4qzBDWRt8mHQq5HqT1orEKMhzotQ/JoqKZ1
5sNMDkC46JeS+THn5oOEcGEK4dTT8E4KbIFSit75/qSIBAUwITuwOMOY5xVJ1pxN+kMoEnGDB2Yv
xtPZjBnOm/Qz1fWLgNf5tel6BZmk9blHzqFC9dfWthjn+dGPl1gWRE9mN7HjAvMzIlpnKnZamMZn
/8mSUDJeRSwriM9ASWuK4vRAp3tDaWwUtebsGdXMj7p90zfsvmAj/xlb2WtNR9LZ7zPI3FzFdP+V
01vR2slXD4xEXyB297mcJDdRdrTHgsPZeaBQDm+my23lmEdFB+N1G1d5bVdRJq/UIg3eQ3cC/L1C
6eeh/6O/4RZgaxwQ/QZaIgq44nKIiLMbeqiZCwJccSTTZ/tuv+nW7zU9pf7AK3cWXm87uswdG8Aq
KlvVODMDp+6FcGeBppsJadhaRlNgzzzGMeM3i4cSLlhEk/ZxiPAzCMWULscXTUuxLdGKIMM3r4+P
BTfWSkJ9cgBbRgDjH2571/f37MSXdg2GpL5+9sy5nhErJ0+D8E93uhNswc6Ps3i7iXMFDEnYt8aU
pz+16GuTHjDGSRMmO5zKzqxml5fwiTis21osjPyi1m7UDSaeRUmRRyDEIOuQzFPEwhUp3q+D5iBf
8sMFYLGhdDQg/II4dhd05nHQuZcz4E5aJirqOQ8dOyMzhmIOguDp9DuWF3wT8zswBnMJQsgy4FoF
J6zGv7KuGipiAv/ox8//JdD27fNNUJB2FJ6AAqwBjcGDKguICosT2WIOs3K4EWvnCpxr6i4/E1pz
lWqnukMALP85gA8sPcU2ykSIZCZHNGDLivgTzZkJ1YgHujHqZ4rDc/+0zDfPSrJdx4eun0VcHDC2
BEOJkrFpwnSmLWdDWshF4IcuY7qDOGJmFiobMy+nt8xcLK/c9mtKRXCpKw50LTmbVhv+8ENaYjzD
AcVkH1FYGoaxkPnhOw29lGEm8Fg03b98sji/NHw8Nou476ZCoOeck1xapxpZagLXQghHnVtnwrSG
4BXYnQiOipaHS6aflSU/lfBOYRboRJFsExUhMdhp1n6uZuBTCNeNXwJWMn9mGBub9qYygo4v9Pzk
Gx5H9rBCCZ1/xFJJJNfjwTP85qhie03WAMpx00vI597ggZvqlWyPs2Tzgvq+Pyuy5ogUzZHqvDpp
S1OvNcI2ZI24NNwsQt04VyVc7CCYad4P+t114xMuJpmDKxt0bfvavVGlS1+YMPJeNxiED8Mpa4Ze
aFGsz+i8QvAYfaH6qyx2z5InEg7TAihE7yYLNTEZwVfZUf83qknL/Zksudgzw8opLaqoLcJIAMde
0lJRcNq+5caS9Dgx76l/keUsIiiopD6TUaldru9D7Gs0h1nPR76lKgw9FZ7WvUJHQDdbNgYXnPqd
HtWiuQLJ9T0zmvTkkTn18arYwVs0O9aaSxSNwEAAZ3QPfUEE6OLRwN5euPwW5fDCJqPdjygm8Qb6
htaks9WhZLGuIUz0fMWspEbYmEOIRhHGzaH8QYjoEd9oCN7R9vELZiQMaiFFgw1rmyiAQ9+utcEa
a/hb4WMADIvcn2qUYCGEmxQCnC6Sf8xq2wPwPQd+rAZjBlmdsgdCzc+P24PWZVNB9QZjI2L7416b
L2bTTFd2DoOy/KUKR56xpQ3qdY/m8QlIYYgkaxanGkf4w6ggkCvho9lRGHnRvk+L4SU6FQvHWRXt
HGIe6c9TwY4dy9IJQgx76swnIsEszgxqyWdDRzsVCuVHmscOnfK7ssNtxfX7NI75xH1ojkSI1YEl
ce8f5LXxgWlbFTV01fL0mi8FcRnyOkcwxrMVvlVR6SFGQmP06HW0pHMYaeVrRxZkfz93rFqaglJO
LWCGK6vVs5PJb+vnO/y74lrRIpWjdYAE4jwnDKCro8vxHB93BrANiwxipikRsgTnpAVlyOzxXtzZ
lCFjZJem/S2L6cEIu8U+KiqDzWx5g+yFFdFFquK5eL9XrUAGHSdmwicXWzj5S7ymzLAn0JLxPCcO
dyhz4/KKQ4TVFHyd5ZTqjfFMvBgswhEYa1hDYyHWM3dD87jzasGSvQfCbgseYZ+Rvt6TVBbvJ+Lh
HRsH3ymcqpeAAUKp6oDb5Ax+GzbXR1IXReIIyVisTshRhRvoK2qyewfM1YOA6Q1oBZSMLLrH5TZ+
9sb6CkGf07N98EyHUa76RxkgQjMsVAN/myEzpeePlPZW63qIqKhUJwSqkJPe82c7F/kFjeKm1+Qo
7LuoADK6GmKN1p+6o0SUnfCnbLZU4JmuvNO2K1IHcT30Rf2I4OhdBD1095xDU6gZmbWuiRWQXHwQ
3vvSqs/6izBn6F7vWUsSQVI1s0ngsKjiLqSd6SWbq0yZEBhNirzMEOMA3PdoTnf5zyvpnld52ugV
Ts54cQmfHyv2NSZpg4b2Xo8qleoc0PIMhRr7SXilkif9b3m8LUvj9NeYNKAEj1CdCnHOcvuQC8zE
fodde6rtEkZjkLAgXynuIQeZltPNGz5HwmHVEzGUzJ4G1tKof/wIlhQHPb0x1YDA9XEVxGiYlRSZ
Uf37anIIJGLx9dXivQx+9i40vfLnV39Vi1pBBNYcBpJ44nQzwwB6E1YJxYMYtvJkwsuVMeq9jxhr
OGTc+irwkyFH/SNdRhOVPisbleMAyIYgidCwOl/Lu9zqWsQJQf2SQXmV91A5RLJ88YLEQvmVOrCK
7XSR6vD6gYV+LGnV0KxFbRqFHRiRVo2U65CjO7ka6IoPnfirJBPl1QuT1HuhDD9DvAnMiOw9OwdE
zzT8lC66SKWuSaHCCvsqAi4sXiStgBMNhUn3lh9DFvIhJtQqARXLOlrHC/GeyOrlaFshOUUxbf98
uJf9zfxmyQoeVunT4+5VPhk09uLAcBoGbiVqXIhD7V8M0Y/bReq+tiisKijlCgtxvj2uR1s8IdCh
wc+t22WiTsiYPiPNIQYKPXd6IhBIlTJvnjLFiPRDdxYV9duVxLq917le33CaVyZ0+P1rtuz28B6l
BMlYpftIz0cFkGjZAc9fLbaxy48/LUCFHSFbw2k6zOtVp7CcsMnY5jPoVylRPgKMeWw0yF/QgiD9
oh2HLqGYEYV3vhj3Mq35AibZyBRl7MRUtvfl72yDWpGmf2+6JHjVdzC60QOFbrNxBM5TLwiiD0Ik
TMRDBnw2WFdEqKlV5FVSCK/AdQR4bhRKyuTuy9MWId8KbQGpp8XT0PA2YDwerR9ikUwGmk9YmYBR
mZ4fmOVe9DHvAWND8ldo1ZF77GVDUTy702kSPICkaCQ8usiVVlSFn1pWNMzVP0mqJdXj8gPxX71U
kSzQ3l/yAT4aPveUxrBxx1RDmTpLQE2alKxB2YBHkW8XIz+wsEPNnApPKpmsYwcg7qYdrOkvWn44
34wGn0otH4CAo3MQCJOTKRjKeHukzM5iccJnVP0YMwr18OLoQvfsrsZmYZn6jg8E6PADwPTZG20l
qVlJocBxhkildoqN5hbqjF4UoHLijOzKHYAYsuXliWX3coWJYp/yD+vWnVjmo2GDRcaBb2WMN9lC
tQ7Y8g7fenr0FvHMbRH88K+cRvmv3ey+bQAts4UbdlyDAD+XSQQibw9NW0JKb6K9i6amUKzRX+5e
AmR9hC6rXYfftcQu0I1RZweKJFD83W6GKFQLtdD0z1uefqF+9b65gBXz49pt3swEev7RXyIYmAV6
k7JkQ2YxRgop71jI/tAERjI+R2caiQY5KbOIaA1AG/Xmx8Xx0gojEBuzUolTiRI9bTvwgqE3eBHA
EABc9VWob8/rvQoMdmTVEOuB2gi+IxYjf1YQmbO+oDIcBySKZUvKbm6uExq6o++T/M+QitIdVM0l
gMMmKdjjCbHdfNHMeWgkf4z+LNA1TSp42S/Ghn1nXxEnxQztioxjfxmVgDQ7LxZf8Xb74Trq5BZx
WJ69nk5iMsbkyaARMNi0zbAEht5JX6PBjHUhZEKctdymLzbxDtIgpWM2xXrHW1ZmKX0bQI/rzvOf
BZdG3mUNx66XPYu3bbP39ik64339xDnLfmMNZLCZE1Qr5m63NoYD2iQzL854xHpZV+cMHWGkplNr
Pb6kMzl7IFnTNIUu49kChu7CWlHCPL9Mnb478UA3j3PgR6/rhBZAoWWDf3fOllvarTCUG05ifDeO
wULjHTUk72BZhWDL/Ge3EuV+Q7pKl3LbaIVPmaQdv/0wmAjflFCdCfN2UY0yX6lIzxIywE7sT2Pe
OLvKihT2UhzT4KFJfVIZqwIX1UKEO7LNIu6nVnk8u7l1yYUZblyNr4ptVoOcSS5qNXeKwtGAQ8LJ
aDNYFAvcIwjYVs8idmhY7aFV82Y5+c9uZDPh9D7S4XGDU8GOtzZOe3lpuS1E3wYc42wSBKMWKsH3
YZTqSPDqsZAatsLGeOJ945lIVp5iVq/MRlGsmXAi/cr0WvUj2KEx8Qk6FsOlPZt+rIz8k80vZVLs
QMBHAcQ0Ow96gc97oEW73yDc9m8gLNA3EFCVfQ1HncDy2+wWYQaqgKg9OYEAJQ63Aq5SG9grcsH4
7wz5nt8Mt8MRdOy11UEyt92NKQvegGhGJTgnUBmVe1R+N03WGH4koiIThePAuzvgiswtvnvt2Z3q
82maRm9YCHaUKNrgpR9rbO8814EUkM9pvlSboN3EI+FxDfwtnFj/7YB7UFn8GqQXapEetGXbbwKe
87fdh4viFe8ThCemJtyd0OTEBXdJjl7E7BX6nfiyP8sVBAnFxoquBNNMEnRON0lzeEAjweicX2C+
Nuc+EawUNx+nDf9hof6sAdqm9VLF3JbI14BB/7d6e9dtrnG8hcvpaHDTUlMjQxfwGzrBQN/g8S1r
/Ye+jOUpQEB8N1oTGalSCglbQcQH66M54NB2h775HnalpxJoxxT27uKZNu+NRzvMD0idK3gS+MNC
2X9mhvCZ4p3pGTFS++hudNQHch/jl9FCss/+jV+HKa4dLK6sLfw5IjNLtu3lqKId3zhG0bV3obM+
98MyKZjjxMTlnYJ7DvssCX/y42cxCHWS9Dn5H0xba6uUeQOiDJ4gtJe/ipKykbehVLO+m1B8WuHx
4BbkZpbr5IA75j+nurvq8g5XHUdM5CUZozDBVmaAgZm4ldn5H7HdwPcljE6u5PPun9gfK3pnV1dx
4npfewhjU8apQW/Y2ud59x1y/jGwjlZIjo6g41+nUtcFx63iHOSy5ajr79cniLVKy5qDyhAhmrq7
/BFDRF3MMmOvSUvXybLmhZZJFv7nazNndO79OXJynf/mDopAq2ZmlaGivmzGelUSVNJYo0RYR1vR
Jr1kJ6cprCkc7kct0itMNFruCZdY3mLMpSifPLWJkq4zAGFed+QYS+mm+2z1lpm4zT5+dezYRGrt
j3TX9K+SG6mxF4Xr9HVoG1I6AdfXu2vz0B6gJhBUcMioL9OPVVeRkKsLgJvUQZMzoo838jjYudF5
vJ6DAvJ3vgx+ZCMpXTqLOHd5YXJMFSK0cc4oP0QvDEq3SmgNzxwYvZHeD7kGtM8sg/gbnZwAxF8b
1soziL3GmO+Xz1y9txX0oVcIlXpKDHHrv4gCzbqpcu2dJAS8HyB5eQGzCefOh6ms0yiXCzhcjGwA
AFrcy8/Ewmq+vdNV4CnD7KoKHuW8Hbj0AZDgv1oyRl8wr0HP4xN6BpUiBXhLzv1xM7zkWDJCivik
J71GqrHJ7EU7+gXqkhMfYbT17fb3nY760Xr5/q/dJ5/jD/yoRhFSHWRQtrCz8Su+E6qjAudvDQRL
YqqAganjGBx1hmTpp2XIDMPCnGaLC3MotwA140G4BHqrDDS9XFN8Re8otvWBFsX+B4+wkU7ldwvk
OD9OVvsrBSyuFGK7/YnbCPuX2HAH0gSSiHdqsajm/BuZHwMmvYjv/07Emc7IxKiH2ly2ptNcQj+K
4gvxzUtB7uWv5XOjAH3bKxu1OG/gOkHI9nk2TWSRaM3U4WZ+ReGB/E0aJqMxH9NzbdeE7OAfUUk8
LJx2xeY56dS+o1QQPATMZ04QcMAascp0ASjdcWguED7+liW1BArLfJLXAvrnm4XxkAswoRDb0kqH
bfANf/BRcJByLzozP2DKbdQVrHxsPNIWRswsNCWRXycdJV8tjJZtBXMZ8aHTsIAytZHbAGClmRIV
TDepiWJng0a7XjkNH5Ij7qb1YYhgD6q5IyJLTcU6ol+aUc9lcM3HJdVGAqKkaKa1TPS/Z1BLTSH/
g7NxdanbdIosDA2WVdkPg7XcI/j7QzYzNSMIG4qKPv9BgIMWMHK+7OXsVfo4oPJw7Uluuoj4Sl+4
i5IlVFEA5NgLOHIJlUvaaplTTNnSY5Hb/Go0s6SqNy6dqjhb09nc2t/7m0D0dQNcwH+vHy62aV47
KObTfta4lX43FqiLpWQjmc9qJvUdelgwAgmhcAISrLaz+LZy8+PjBT+IfYn/SsQHhulnAB8o9BFM
ID1clJGOHVRb/IX66nSYNCZp9eDYBjRNP8U6bvybqVWgELj6UxFb0tyvX/a1ixHrDrlapcF6uXi3
KD+q20axRKfJ9M/R2egk/V1fjB6bNq9nqLSiAw2cujgrQaRVcCs/UHekLSPPjMhLGw84X5p6d0zX
fpyknVHG6qzs5rV1L8q9EHdMfPYdZApMUi2Le9vyp1K8Kqj3bVPX0L29z9+w3zpIagCGWp+m7uSJ
IKYi/cqHoJ8XNix+0L9pibB+KUK1MlyEPj1LpdY/DfS8WidCfIloZ7wTHwgIAXKVO68siYwe+Tyz
yc252oSG5+SVQE4+ALEhcA8YNQZqm6UyeoQN90ytn/y+IlWR26PyQO3ttQWjR4HMUgxnU2ObnVti
8yqaXpjsQjf0qEdpvEz4Ah7AEVl15RuRQXM38IVzyAtNQyJIqSdp/IVyJ881hzk1sM3u9ui9vcbD
NrebiSZpVTu9mFhKD1R1AhMSXbmdCwczWaw+r74kY8eF1JanjWZ7YX358N8KVC6/zdM8hNdV2k4N
5Ha0wraXcQXnUcE+82SowZ46HuILApaz02/LPaJtaaEuq9/FZdPpAaSZ/aTixfI7TjRya8sAMSVj
T40UCGSH1yVrYkDjq1oHsAQMW3CL5/+oaXVkgz/cP+Nlwx9CUsKBD5cHCGyAzv4b0AAg/dPMY99n
O3xllDQtRCYHvXVDMdhZJEAQ4/2nXexEraDQualYoJyI+yioQFpJSuFYzKIYApFPuVbeWiXfn5bU
Dn+og128okzHCZBzpi2WN3LkOeVLpyZkVZwAS6Z3ugw6VUmWySr2T8c9sGWZAjpCC8m7+lcuPTxm
dm0csec3v4/PzwBWFqXSlXbwYlWiVZ0wKyOr84i5lAyGm61z2o/pCDMk8pM9JVIhzmhNpF7DoTpO
8Tmnp6qi/+Ll6KZqA5JKNPeqIUJ6NRHceX1/sjcZ21+2sRrxGSrm3FDr0FZbN+TgHnsWFflMssn1
ufT+uS9srsMQ/u72xz635LIwO7EUJyrJkwog0h36vMsNQJW1s6nxRP4TX1a7QP+3C/uXoNvpmsVS
xhSVhjJU6/uCm2AtYLnAYu4ABqzi+2DD7xROfA1g2pXpgvQPqVeBxJmWJXfwyEAlqQ4Y4s+y9ebn
4uucOWluYC89VtStLQ8QCobBJZBcYxOSZrALIkU7/ZrN811Aw+AdTGAW8W9hfzULatR7WELnirC2
g4++tdXAxS63lu7rtfFRcNwxfwDnb9Hk8Jra7ZvKN48eBlDUWyXH7/tlsb13ArNTWP9MFGAnW89c
HdEMjxH6PtM3hoa3QY94irdtue4rydDXz7dt45P3nmCAKLWEIlyRucOaxKAv+2uv9WzkohykxS2X
eTeW1LkCwBv31QI7lWm1WZMcVIqI57JJxlQXBFMX1RalbE/6K/0HMJ/+ePU+ZMUtRVyfQr0v4Fd5
iFJ1MmgbvneA33ZbLZC0meUFRq2QYCzRNZVD4vpOMl2SR7oqvhhTqQTzxTl521DzBsRDpS6KMDTd
4aDeoIMtlwbhn9hyV8xa25f4N88I6a42h+7pxMp039K4h5nwwgFUskfmLR4/CN0Aj3vZL3yumH8O
fZg6VLPD3ZHOhQU8RQB7YrOkttKTLUSt5OdRrOe+4xTqjXNcNWuCQPGXdkRRuKKFe+tdddqAjTLX
qu1HKVFT7Ze6Vdgy3VH8Fe6+zB55oU6XYaMh0p8ygmX1ATQUeWSm94LmXvNHU4xuJxR57YBVnUCp
N2X7S3rG+famF0TgHhrRexjKekMQQANnJUcBQCwg9XZgXd7BuWzzt2JjZCWV3JtmOo1R8CFeYNWk
FydLo0ASVL7zx9ieFpzF3NiHw1cVu7JZJnnk/BdDXi/U55/JaiMxzzxjo9E+JJ9DQxHJP3ZnDA1L
GA6D5mZ1OKUAW19LMpoeWLmzCoeCFTWl+ZCg8Ls0V+TxWOTrsiGxKrsMGGQtJNFviCKau3gDOkDs
9YdnSS9ICfwTdObFLfq426BwAhMjWaXipvlEJRTbvd8QkxNM+BwuDEbhwUGNI0PT8glt6KPmR4E0
UUE5x9rvoCa0Wh1cg3ZbS8qIszgUW3363RkS0Fl0jZhIz9VY1CMiDjb+MCFzdrUSoAT8xRoTPOBi
iwo5x5c+SPi4v8sYn87fzzYGutZQTgadHZ+OchXXLIG+7segH+goWwQEEVlbLVOBEz73DpLRLuQG
AwVEx8qkCF0eeNPk5tM6hRA6boaEgz2/q3zHcrTRoWe+d9+XAhP28lhDCmNYhIXa4U0A/I4h4dGZ
qHtvjbCwqxANu0APk5H708L7cLdTv8jTZFZtJXtQBso8iZKGri90ant7SNBBVSUjRd8PxyAzFpxN
OgnXPgRl9EVjVsmVt/2OxONGxwX/h2Zx6B0Lcunr8v8se7nuQGqfIC+YTnGtYZytg+CbDBnTBlk0
qyawZeWEEoh6+XfnA/0kAbnTbiAjtueKNABeRcPgGBSI5682y0slkF0xjnnjRSMfN1lfvtrFOrG0
5GQI2H12gu+6g99Zb+WDE7fyVM56tBnIFhDBkKItcP81HiNKAhkhdP5BBuodlzzvZQG4FrSbpG8x
8iXYRL3LrftJdhR0z8O10OolTERdUx5s/l63qjPKgKwoegRko6fbEzuKUAtG3Tqp5Q5mSq4RzaVQ
xUe31hrA3Xb11471T1PTwayko4AsVW71mBGesUsp3CY2WiwvMJPYRAccNKcYfJkS2W7Ie0wwCKYD
+TbytLVJPN/fG8ZFXr/G7yelgXbjpSbBJOnHvzUi0HALJBN6PbQi1Bh3iq+ou/XSJcqOLtEpaRs7
zDIDT8Hg5sVn46Nl5kVkTWT7P/gCMVcvdEPzT5pX7GShwpvTwHZAtpVb6NKxkAJZqWsrMH3jjoxN
4AGh5mwj6As2vEDWn4mgOQlPhw+ors2XyCV/CvuQ15D+oGi/q/AGczx4or+Dbw4F5OLUewual6XH
pmNv+21D7ed92GXC92aMEuwCi/tzFuuTHBNi5kUp7UBP18KzyTL5nrpE9NVvERVhfMBrTrbrnr+O
nKJedSGxUpVcUt2Ug0EQh/KC7MXuNZCZdM1W9Hv4+80ooYQK70i2bgJ7bRbT5OI/0e9uwsGiU2TC
eOmMmD2dJvdhXXDfxebGZHND0O90r9z9NU4NvzRvJ7AVrt6EOwxh9IOxCiK9ix08VsH2DtPiKmYP
bGm0qHmR+wV6ID9UzqYU4tTc3b8b1cs0mL2Cn1l7vXxKVGdSdCpSvS9L3fccTGFk1K9rauo+zofs
/dgz19iv71fi2lL/AMvF/jEHKd2eMJgPXPb98D0+a+gnQcLTl8oONfiav3s9oHFaxVAsZbbmRawW
L1kQG7QnpMbXW4lUMsEeHf4ioKtEkJ1NJ4f9IVjnmsecSvjVzKYtJgXeGfp88CwsQqrhtVgUiKeQ
F9Rvas/RYkxTDHw0SxI3JWBnqZJks/qd/dv6CtNmQWyqdwNG4ZF2+e8Hc5hysEdBjqRdhAQpAOIg
1tgaOetocxl7BGJb08woMdFxXjgWMiMP/P6dFbxWpQ+vV2Wf2wMMObY8CGV4JRQ2opY/cFCKQkXI
lQ+1kR1UmxdUCR7rQ+hjKVtJQrk5B3IQFKO5gb2b0scDehlNRIF3Rg4qEcQaAYkd3YymNmlG+7L3
Ew3khm4n2ZUKZz+qJuVX7Z+A/8YyQTb6X/7L/QSfJmt8GK0V+/zumI1fMLpTzLCqErqC0vRGlHR+
oax8FiTL55x51FoU3tttA+RnMm0SYkn6sSK0meOvJW+94kFhMaLxVziDRTp0dKTlt1lnLms6okfX
tWbNTE9Q4FuOJAHR3x3WaVF2S+lPL2hgDmV2IJ/d9Q09kRPej0iSBiiO0s8nA5g8Ps3cOWHO79Gc
/pM1rXinm9TUvY/V5F2sS2OpLkZoledZqsYXd3VjwQjy50rwcalu+lSDyVL4Nxn1+GWtndEFDy2Z
Qc5P4aCvd6EKVa2ef4Dbp8uNhbLhnogSHIyzqCffSnqsnXHuqaSfw8mRxDN2OrCEYm7cp7M9DpJQ
SSKiX2INm5U0b5mEvzCTF9S5Idss7RDxjgblo+mkPxwL3bQ2y+nLLGGFMxWJC7oqFcKeGURtYPzZ
WmuLivbWytAg3W7qr/KjJRGFjcdZvugpGziDfV56thtvMcX1wfxsuFjDQn7HPyOMn8X0C09UGJI7
4/Pn+oJcXzHrw+qe5SLEiTQ6HqyslGycJ+ZeaQfyTXDSTDSEJgO9zkFaKZW7rJxZs6JKPJsKTGkw
hgaJE6BeeJCzBZlzZeQd6bo2apfqmk1MFx1blkK9WVWvgJhaOt8mph7fJZVlcNqMhy2EtYCHmge0
M5jXd2XDQ4DW1WOqABVAvnRQhBbIxfB1809VIrByFRQW0p44hsGn1FyvhQL5ZK6Ux2Z1aRXMvWhR
mIFJ6gN1ngp6UZfG0sMNTwUTRq2d44UFewXTObg5KsY8S0kjOz4jJt3Ah9PZuqjmDCTtWbHeES5D
/McoynBJd3w+NB381rQPjH2NXRLPLZU4IOTO+OoQbJiYBbZ+cXYZ7yayZrSDxUYn3T71YiNOKGKQ
594aWTo7+NlDkusXblzUeU2OfeABimqI6S8tb8c4E9Q8KHYO/Bh7/ppuGwY/Gl9uY071tXCoGsP3
+9pj+VCV5xp+FYUv2acl8yiYdojM7f/a9QgXFM1Ktkj3/EXNa9+e2sGwnuN128npr4+dPJ0IPt+Y
+/gr2BS2GKOSs9wZWz7ESVRqpms4rqkpAb6DI7wPY86MLikOFZUzOzo21enwqVhY/YTe8FcBa0eY
9qzYDRAs4nK8y1wrbCdqR7Ydm92VX0TBPP2rRkDysyvKTC8Fa1h4HA2efrTba67oIdAJkMAZpveb
pwoq3GpwnggBLbL1CnZkvXqHJK/ZhBYPgeyvq6I7cv9WhYLWWqDsesPDn5MI12VObkUSszGhDZP0
mY92RDrYIKjmHgPAmQHr1klIy5ZfZzrT7bK/aGe9jftpjcbRCNnqZ90A0yAnj1aIeddKtEiL/Tm1
QqWqWXa4XhqIRRaNQ7pN0i7i8RkWvtnYGgknH3RWOMRw/K5MaQaQQ5y0BS2Bk2TL7gdAt5vQ1irm
ivTDnI4afjnmBWaLzATcdZZTWoG6wA5360PoB2lg/WnkUxe2SBu/Y4EFRO00Qd0Jx9hEXsIipNSO
DmJSX/uOg7T+slt1AoRo7QvDZ8k+7zLm9k3oPTaQO+Ks6pVkboxZPsKN/eXoUK7bNPjsAWtXInRH
UdTr8BDCiN4CxqV37kOzEwkqeuubbhI6268VE4KHGlSBD8Rxpd+1peAxApArUBioeiIMI3EF96FE
2nqkzALcySLfPcrk4fYgBAAqRJ1t/4tXF775XOlcMqaMsG+7eLARbm/TrjY5Y+dcdPB+4e+EpaDW
QzSc199hd/K5ZZft2UJMrb+mNCuQxCgOuN7puo2agcY+HrRgiOp1RNwcGFA1FsxAlIfah8AV4Gr1
ks6BJBLhX62PqYVp2+8h0/frKt/2WkBP64jiCuiUodfsvwpTmLDJGi6Cy9qm2iyNClOVpRRrv8pV
Cy/ZapeOBocPIzhXg8hKseoAwB+KI5qaPt1Jj0Gw1xV899yG7fhNS7hBAzLn00lIgQ6sNbmKcRdr
c/TLeisU4PhYC2NYmUrIMvVTA+1fqyp6roQ7PVoIss/M/RAgKBiftM9p60MK9/VWlxUsAoYvTkrA
/qtSDCno2OPOM8/a67XaH4Z2c8LdZFghGap4azOvOgdFonPS0H81O+johc3Yz6ViICCLnRne/8nz
np2wW/MMAdc6Vao+M1qf/CNqAywUzGK7YUI9wkPGcGGU/PwHLrh1SS7Jl6bJISbjXniJcDM5JmJC
0pKf2v2f9RL1XpZ915Bv1n+Zd24GzYlxpx/4tsFCFhLDGo619jQ4jeTBMIK0ZbwYpKGqZytSvRcv
a/r9yBRN6t77lef5kBNgUcZyEJEAGdNUog0KNKZWj7JTwMqg1yzeYp4t9RDS2aOOV2R/QRZybqL4
HTUuXbpeylfPUR1dHitApx2xrDc68Unv4+lxwafJXZJsoAV4MH2fz9lopR8GMtz+XG+kn7ub8IlR
h83Ckt45l2X0AtqjfpEZlDbdKzmW+1SkWAY1dwidEG3c2GlDrfQxrPJSAAdJBKjahxcYy7VfIMD/
5q5r1ZHiF1fkcPhDzB4Qr9jcISugugLwTAWyYU4MZvHyLsfOt4JJh4Cns4rALsYuKca2G6+Jv/6F
VEs6qPwr6U5S+4JMuM8rectCTKy3tc9Rf87XeswWYhT2rrYCaj7d2CWtgL7g8uVgflpDP+uiKSyf
Lp9YtURai1W3KFjszRrdUY+9KGlRkf8tBtwd7A5Ruhay9o/KFrszmhfaznXmH1UEUZeVI6KTG9bQ
rWjUYXp3JVvEYGapcWwDlQmtkA8ZD3tlp2KbyhoWrB/BbORiCTPQlO95Jrh8T+QvauA20Dd6Wgzd
X+PSgjQxtPbqao64TS/w+NJWmfpYcZFCF7PtCdrwy/lc/ptoDf6kGcq01ZnOIy0c4DAJQzpwQVhW
EZh6RJElfuH+boBP9rY7yBueuXOEsphpsciYzDq/+rFEkDjk3YwmZMryBmmKCcepwYKWadGa03fc
X5PGsKIq65rdq98KVZDzaZgoVYAz1euDe6IZ6tpTyiiOzKIEtGwGRtysPgJcpW5+s4JLLgPsTKf8
OluFXmsx5WqEdJ8RhrteQoPTO6zDZ2w2dXpXBXytBHQ8IzIvf2kcSnlOyAxdwofbUYOlksJtoSRo
py9D7ILFN8Hqd5lZ+pNgzE4KMOJKaT/QW1p0ZuRPLgU3V+JE4b78KR1FqQo8ZnNXuS1kbWax0RZC
qhm0IW5EnZLdI13Romwdqw6cJPBl0Wb5gd662CWlyzWIMyVxmdI57nNqMI4vJ1+V/CVD3vaI29S1
vkPbUVneK+TPko05cqP+pynfaknBSGZzBKWouPYhe7e4KUIbiKWP2Ovev72DbHssV9D+9lUJMa1F
sWS0Dcg6W6QmfYINjEFpSwxgBiikSLGhx72dN6lYuvKrva0L9PNitkCu9iQlSuaq2/PKcJmYHb1t
GqmcWwTrT+WEjZz9jLreK0g1zuHFWo6jU3yTNq2mvYxQoObCi5FRUtEnXhWpT/6KQ5P9VRyXYRIH
CYW9CgKt0b/XzcUi5POmT6ONdxOIkByqVUWWxHgmSRCzql9lQmjsOgrTahjOz9DPROYqKNYpKZI7
iRUafNYKbIq9fQ8ZEAk2VNN4XbedAIC4t4CqImI0okpnyZ12vwHR3xLe5uZ8Z8RH6Zsngj2+efTp
WhR3taok3hjHNyUq5cj0igxObzNX0z/rDSdXBG6gpZC576XkIJOjyhMOBaEaKgAdNMiLpA/LwufN
6ly7YBJEphajTPwIqq5Ez6wzTWIwrkDK1FydHMK/nnqMACzvqlMb1Xiell12AqKDtxes2NzGXth9
PFCoTavINFhGHNXkkCSU5zjVDiOh9moJNRBa48jz2ONITe20/WOh1DC4ogT48jmFOsVHeYU3bt3w
zhB/i2btZgNjcyUfbE0n4JK06MluXbNcBLytg0REOs9wg93NDNvRRmbK/W/6bBwpdng1oUHMtyjM
TyBUi3vvfXFpXUKzO6zQF0kLmvb80Hyn7jJMriGY/kni93tVZFBWlAwqiNyL4ZUQUXFKlWlH7853
Dpfo+XJ/yiSWQiAKRIKNXRfcLR1nXeSKG0eaxFWmuHBLURe0po5uFHH1fIf93pFSh4yzJAMWDV7y
c8zmFShNuHWuyau+6zxCotBXfP+lFQYfw9NK4wAwc3p8imvFoHlaMMuPnrChqyB21rci3rIg4BJQ
mGkbcp/A9qWOW19EKTCp/VTd2nsIdoL/L8x3IRI2jSxr7PhWdM+fM/Aahx8sE3yLbuelsk0vTEdh
DyKSlTeQnpXQp1J4lNUqecmWPw6LQ5qoPQ1vTOpRMzV1suagvULMWuoJuec6DcY1ZWtBVh6C4qFX
U0FCyeGG0YeG49gIHOIAYHVT8nkf+IczZCMyI3ThOCbzSK9VnkraQ1Uc9THDIGWbgPpaijqyVhNH
BMJpVfCNAGX5PTmyn0jdLEnL6j0W2fCmwUyLDJRvIOYm9E0VfCfv2EAxyOpsW9KGii96tpBfLBIf
q2xnD000ncmps2k5DhJ9JvbwxGLwsWUPdKhaE1XdV8i8lQqMoXxq/fh55dCWhmXrORXtZL+InswK
e8g8wX7LJ0Q6x5yS3P5QI6zYy62FQda9+SjPs6HV+R44DhKlAUeGOks0qg/ikqu1MzxQDs1hdK6r
7bVVh5orvIeNBCuezpGWvslRzXr7ok89r9qpboxgvOcwMPCQvZvkOEZM1JgtO74LXlluINYef9hE
v6GHjsiJrfKfI/KGG+LluELGpNrPq+HoD9VZYJ19/iorxJktd4+MdTvxX9elsm5RXMzZKhW1oZb1
L9pYti0w77yEukplawpgOm0zarEV8BSP4pmo/0/ydF0YSfjZrGUvruyR68dJ4AQkR6i1lO0kmz53
b4q3fnlm9BN2z8tghAgA6HOIz39KsQqHBKUIptvco8p7K9SkOHQIv4086pRE1yRDwDuxsnBL0RbV
S5gA4kRPmUXcthR+ZS42q/qq3gjBMZ5W6RFBRxrPEP+3pMeVOYn+BQs/iwQT3AjTEcP6XOcssFfC
8lx9ibXiE4jjmf4ETT3tr4mtRnSXQvkL8iO2ZGOuZltPP2/sGXrhImEioMgZaYVuo48rksrhxt5h
F8jK+IFoSan0OjjEZlk/AiZknPGvyg4RCKQ8Bb48JUKnoM9xzcD9JgCHx8I/GDofcmV7JVJRfDM4
Cxdfxo3Dr/8sSyVu2faFQWjeJiMWnNy/NrRI+qdY6tlzyT3ZafHXiXq51tCKqYUWZk4Pqjxs/wVb
+nw4+wDQWxbXxgEMRlgGZsjoYy1UCeKA74UvYBlfAD/E3rTn6LLs8ncLLvVNk9CZFUqWp8JuUBrm
GfbLpRGMbIYEDdJ2N6Jblozp64tIlYHNQBbDPfyOszszWpsX9g2C5nh02oR3ONVtxdg1cQMv7m+G
BiqQXrcTEptJfl/Dfr4ZW3garXzJO7OOB4YgCJOJZy+YTfzvUZhneD+fmFA3N7KZjntIt+xneSAX
HQSR7PgPo7haSr6/fN0QzJlneLAS+frtUlY4+iwDRpSCgUQYftzXOXi2s3+pGs1lYiFW7M4m4k7f
hu1kMrmpYcWvh5PQz8oWP5SshhAHcVHgnfLYzj+k3W/WAc4OvdmBD/9+2fJcr4G67/sHFYhvzymM
+oYyGlRvms+Ks08yaimf5pnOf9QzNhEBzdgWbIgSadoAff+Ty9foX43GtAafCYeYxhZpegYYHWtQ
UYliXnDRafLXb78bKFjhvUUHhV4qR31Acrq1j02cQm5fhmOjzDZNnu6ExtlwXLiHvcQokc7ghYdK
BgDfdQ58gOaIvD3XgVlqNoMBHtjZTvkmumR0jcr5k9vsXxwRCReH/+Sm+0G2LACHAw7uVwVh/hXa
aHDrE8wZR74wegq9Vrc9Hw/RQxdPFC+VlpWtQffoMK1uSUae86fjrau6LZBd8XS4GyQHjVLhsbqg
oWVbdF2tpHGecb2JoZlJ85EBh2mq3lWnR9Kd4YQFSMnSTN8NqrIFpJPokRQXQO06pJEWosjUSGed
vmiJGn6EN5KO7oEXFcG+zTCIYZkN3MFyp8P79wNpt87QJhHuMXigNcy1OFqP0vl3+5CgJSDe8QpL
meJlxRzL/l+bnsPUDzZ6Vxl1NTlJHeynlHZg6K2mGDZQ0/bed2Mdg9YA5Vazir+VtbGZsvlTxE45
VlFEy5BlvXAShcV9zYpAyb8pxnpnlMUZNLgruE0pla8L4ILrXR/Yg7rXsg+0XoWFOS0jZX7ieCY2
QX2n5ku8MSdA9s4fvgZ2r/nqbRuhypQtAO599kViXsIg4aR6YVROpZFUE65OzyrExSX42ZDxSHPI
FMHhM+3kkKwnWBEVjmd8TjTlp4phbVnB9LS0CV+B0jNDKwcjh5Wa+JQAL75JCaDQ9CzCP9TnHgYU
0HoY8DByBuAuUHPOOoYEcR1f3GK/mSPWu5dZIRMGv96GgEUbWEpRi0V34tnR4sg5DHTcSc2tFWmB
+X833wwCqPgQwV+nCWHpefqRiJwP5Sa5a+l/zcuRpal+iKmMEjOk2bh9BpjhPo0SclJK58El5JiR
bWk//AB2/1jtiMkhdHOOiSS354pPtTbdBBeJXwy5N6x1Tg4RvjrTj7Ls2HmF+UV5kXOCSJ9Gctz7
3Xp8WWb12T6YVskpV/xOCWsiWa9/WcOQP6W2E4PlpgHXN0GBTsQghYLueK3fVnX+U2f7hI1KooRK
tmddnsWtw0PRj93KDQnAnVNQEzkJhC3ZawxxbBcLQVPv6/TBgskESLm+voKt9v+ifYVZT6kn+ju4
VnQ/LPeJ+3R2euzktVNFAyKFE3yqfqOdx5JqhwP5f2qpFc+yN64ezPXVfXZ5KzYbXaz8omsvFH6O
krphvor0jCTzoYpdgVvnPP5U7ltOwRho67zl+DgtFi79cBTsJX7eg5vqi404+8xUiMFoVYDoAEaL
+Aj9bOWQTDZisqtpBJcOlvu7ppQUU3s+CVc1VIgDpq2ZDxhMSbPamN6CKqTVcE+YezNzrTJsVl64
/f9YMmL+OJ3Zh4OzYWHI4ISDE5ziN8piI3v1iExvYUBfoN06kYiCSWMWxZ+opkfSDHhV+0upxV1P
i1gbptCs90UYTHnxyuabznajMRXhLi4E3Q/l99TLwh6USUHD6RIErklHHjnybzdbdG9k1AfL5owr
/k69oTD8V3r1Kqew8dHqD9umqx5IO8oDO8MHt2arusV1qLKk12STMksl2quqc+acDjtXdDprSSzu
UDYWIXRTJDuzCn+murC4Kd2CS868jK+BvphJ/X2iS/zquOoiJOFbRmXeFpBFLGdxlcKkVbr/r4Fv
orshlzKgML6nioTSRhdUQYnALmuCXXnkvG/EZHschTGwENa1uN367EfByjh7uSUN5Q4VEqZxsrpa
disSswhW1PqVUU92iO/sa8f0hMD1JE6Rb6UEAf3hCE9zAzaHncLebRWwgb3mfS5o0N3F/ebSLTiJ
9PNHgGY90+QdRtofKiEJ1arbzu1knYQtgTlKCuUS1I+Qs+bdbyA80PytuXfZBh6vxCfhmascRyig
Deu4if+hpZmtUY4BFC7lenmY31Nle54x2v7YeW515Ulkrsctp08F3nr34sU3xYR7oCu1XhRRZcc+
W2bBpZsBse93eLlP8M4jSuGZw3C1ARQbW6VODDa0tZTCiBonT/41xyxO+I2eKgQ2M3rIiVD/yRgk
AI4BZ5y82tQyFzzVgOo+MZzku+vTgSL4RpzCV3uWin04vevsf8KUzRreW5o90UONuBehBJKCWWjs
A4Gbx4DxeSFmyguJ4C09IYtpJijNd3o1qZ6v5HKJPhhPfm9MjBpttXl4P76b42YmD1B9hMbY0I07
zu1k2tUiErGHsS79W9vH1Bfox5ywiu7fOpz9LTbq+Z7IpU68o6bYF1Tjo6RvULbtSL6hUvNhTE7S
JKYMNU3PLWtYd/RLwqHYF212W8Qbctm0jW+HvcaqI4v0RiETWGiD8Ar/ZR2EQAINRtHY9XWmFa3h
47X0k129t58/2uxBDy3PWVxebT3+Vjk4OGcyinXsItZmpm+29V7zVhwAPDvcVFLiZLBbnGc6lGwe
THbRiDyZuCzmMIHVu9m95igdyIsdWNuJ9ixFwfFGdDIJRIYLBiXPD3/SFqdGhPJvNydaua+oucWi
J15pL9V+g0GLto7jc6xV/xE46rnd9c0fsWbAIt69gqRMg627P9X3atbvvva1QRjnaQA+SwYVXJPp
ere+RfLNtWbtQsPtRSPa/DJdQqSNN0zkjeFkq48nfNFAr/3XpY6znN3T9hHWA/KNbZHCuVwlm2gF
N4BJPYtEe+Y18Wazb9drK727hdZQ24S5DOzFFBxm/kGApLGjenebR/B0k/xMii92Od8XL5i33n2W
jhHJBGwnGLN5O0TGfS5xAMWPR3sQcXOLZAs0vKz/GSzLNxuYqNnKzvQAeDzpfEsT+1utHBC7GSBG
6zRUFOoTsfKH60OzMwndCUh6XJc/wY+fGBWYUMbXydVUxeNe1SBt9/1kpP+k5iXsh7R7iVZVyIBh
OVW2yHdubzvGt+AThaHZFeZb6J//f9ZTZ/zrc3xtFaXwh0s3UYSoL7xu9QzGaNaEa+Oyxi+29B7P
h9P52dE/qb0TuSrKrFy+cLQDvkbhOmJr/JIpKczS+rkBdaKOiq4z5/SauNR8aeDb+JXt8tCWV0q7
QGUg+TZ7VHlH39kPc6rcTqkdsPVS1LgeC3KK9FIbE+0QWrSZ90ClAkaXEk/wjkUZ3gMWXyLyllEm
tkEumgKE/tlhg4eX/ceX07Ug92933zNE2yx/bKwt1AvIiRVm6l9hb12qX+g/cY/N4p4U2Td/QM/5
7UrsvQU80xgKcKRUN65jaR6tM5CST5qHnU/lxgp0S5tMnIN15B8mCVl3gvj3CxlzGHLdKsBcVBli
wW79tfM+71KFGqAsmTbQ+yWvgzmQ/546iHCon4FclFXHYYu5Ied6SKNzGXAP2jXmADpvehUtg77y
rUdXGofWZRnNMb6Nhhir31pO8oEm4qjnnPX2jDWBswbCffTCsAoNkHsOXMI+7VtTMlEr8M/u+BvT
1t1IZKa2JYQ+zsVRprHlxAw5YeDEKTmbyMurh8aJSWcIIvV9bG4JMpQvNZUAvdp8xV77qBD0SNID
+fCSnaWhMDUaGBCYqwlkuoMqpROcsIbTiR6yI4V8LZ02qVzhdI1/0JVBlNCb/urH4Xb42CXHDToQ
cbPSb0SmeFiEfmYSHx6snoL7KHfNt21eZoxs9EtTQwbovYmia+DxkOQ/QtZ+PwprcOxSOCIAC4cA
Btcy6hZqKjbMAi5lVctv+sQU4bJnW3sKXizHmRla+AHJD/iETyxAtq3GJqkhYx9deZPUGhhVcObE
BEXB273ohBiqfY6DEN5EcueiARD28SGOC0pCw+m4J07h/QPO4rJazrmV8gNljKWLBfh03PjNcXCh
liVShBL3IfobzEeb5r5L5pQwrNYzX3XPjYQE+E0Tdw2EcPW5F6S4SAZ8f83YKx0qZ+t++VYIRLYp
6uFOGag/DQ1RwqVFZqNAuW8wJ+5nQOa+M3CUrdNhfXWr3N3MPSJQ6BulzRiCOgo6yfDhkKe9i3IK
NH1UPBaAYWhi480UlwLCwduhm+NtuE9Hgb9CXpQXAg69L+0l/LulZbLyTzB88rqer2A6abncUjDm
3FmtykJlCn4kbSaQLf68T7q7iKSEdR/TTU70J1YvFf+4gVu7qqUhUBhQUU1eldBP+zQ9cnO/Azxl
lFfn+Ybr9+92Xq0hR3o7nJOMsVQJX7qAPT/QF58qAs9TO+qT8BbVqKgwi6DIs189yIidB5AnqFWP
GbXx1aU0w70RQLL/ISeKJtsL3H148Chxgv6do6WXxq5HkpuX1s+tPEipo1HSVsL6tmCDfXjV3+bd
h4A9X1ISCvegnkmJGNATPKxdDBcFRaDoOT6OsK4d9ianSuFp9jIm8F2AEhmcSiaPaq+JdOdq416H
V3GrGF0tb3s1bF06NmD6YOMDJDdheGTCQJBVTQSWz8qka7OsAocTV8mllc4zMYXxfAZ1HQC/lint
4hpMhENsOQwUi6NiLca6US8De/vP9QM00ps6b3/1Lr+o+PSO8ZyNr6E31IsH93zOpO4yc3j9aHN1
xdeZa5DZIDwrJysXaEeDG5sjulbOJJzs/kZnVu/HpnlckjRnFJNuf8TKjvHTUBD9qfkoSTeXoWBB
f0MqmOk7uxvopkmwCdZKNV+K8eEw/brk9hNgHmy+iEtMiz9S+3tn/r33KAPQp4+NHtsUHfsM+S/M
FkRBuxTXHFwnXYkyP+aEziYNX8K9x3DQPTH9jmCOy/YaWcWCaW7s6OlYF7TBT0x4JYbV7tFO7SGe
TPx3K+0ZOALSWonDp1dUqnzBZqTdnPiWs8m9mBhf/B/lG07+4B0CkZYtHgMG7ShPlRsyyrKrRzO+
L7dxeo+uFOFIuT276hqqtyaWKl9bcANewDegsUYuhm+w7KKjABPLQQDQAHxJf8owaJaEYVUAWiv9
dE3Mh6N/azahzoA0w7SkSK19i1khnjWYBSnevk73UWCJrQHsBeoRiwQ0i6MGnF9LOlC3OkNzB093
pRWAxDT8JwJl/s5PXl7MqZMUTAXaJ6hXHWHhf2DcqJ6JI/M5lS/o2Tx/kwbFqlSAdWk5BEy0irVi
mO/xAWN5Jj+FIO9BuFq9GSn2hLDzi5IQAEK006ndQw9jGXaiIjQkF9jQBw04tknJuRirS3N/tWjz
s8tFYIUchS/ZBfguFEVALsvkrMjIPl5qXj8X9aK+qS0tegSvS+ZX09bpIRQCGl68RI5gVbP/eHVD
nlyjE07703LMZIfMN7/ONkLNOqSyWEeG3ky9ZktU+sIkAammCEXUhQCBNurBlQeKfiSWgd3piud6
MfqmAFX75atBjZcpFyfIN10pBejYzZUMIVuQx0fqFiLmAvRQl7lG23RrpRzoldiz+0zs4Q7o3RUI
HnzAkRe6NL4IP6JumAd17kIj3EydBt0TWSto0n7jWMzPIaUg1OYsHmDkVkpWCdyeVlgvG1ISHXTJ
n9RP/PCNozX1HWQpDNnNND0UqGrgsE2sT5hO+WeFpFQlX93vc6NO0DpgTweN0s4d2x8KpkRKdeqI
3hK89HgMWqlJ1/svlVEKVoJFZBp8ZTbCpWVfyfT4x+Zl7MGIJu5g+bwkHWQF17GweWnUTTWYS8AF
zpNNaAztVlhHaoj5yh40kym2iYtv7orXQG5UuwAamhn9k1v4WzkTe8YZ5xzIdaQxkTfb6XSyw45L
8kl88yYxMJu/WjruHPqXJtRV1ErTc3HZ7DYYZqAevEePS+S7TckN4ltZfn3UnJDSF2EacL/o/sgW
SNp86tV/px67PMXnAbjVeI8yev/q/4GTfRr97p+hbsdW0uzfgrhW4GHj4Qn7Hi5pLVaN520Ai6Y3
gguoMEiVLKzSt2Ipz0ptciuByZdhrlzh6GlzPlNG4OMoiXLxIPh7WjJUafsSrXmIFdJ7HqhNN3l6
9x+Ip6GId1ohtR4KbceqLIZL0+vLPcJBW11WwuUGCSc5YPJwe7MNevp/JJY6RFeYyIfpjjDbWZC3
FYPAzYPa90o93+vPy6yEVq6yJ5nVLocQZuDtAdlnCgAGBChaA2zbdPZykzQKqoNF7yLkd0NcjyE1
ZUNHEXtOWQkfNKmtTjr1/HL43sgaPirntAtRfl+Wu1ygV49hyRMhMJVkq7Zx+G97fTThWbhX9odL
6QZVnL2SXWibmVO22d0g0jj42i0YCzoNuGuGBOJXf908cOTtsxJXvCiH+v3+kNjQOdBudLVSAT/x
FcEfCuRNCELNbT9vp1Hdrh+NwjR9WqCERP1oHw+dbHWy6Wt39sWvjXFxl3t6xDMpedcqp62hd21T
xX4FrBYaFItV0+bEh8uwiyk0TKsfQUewpuWYMGootRYXz0a0ZWr9fv8kUSnGHfVOzjitJ9pBE3KU
0JzeHUCO6MKrp7oNb/AmyoSUY3/3AtYjccM9CSPpPJHBPZjZYbKdUqbrJQXCD7ybvFUBzhcnW0j0
EMWaq1Y0dOj7CIl/ecmjaJUV84neBiSnZz4YsRs3nwEc7i8t01DvZdjYdkPXKKCEZW3Nd6hMgTGk
UGH0rHzk3HMM6xfIMQQtjxxM2CmNQF/2rknp6rRAuAQK9m4XVQxwiv8b/JMChtslozovhov4M/xz
u/aIymFj/o++OSOmSd0qqCG2D4eZIplkU5ep9BV5J6GE4F6dyMJyl6PV5RDhK39/GTucdpobmCDA
om5E/NmfzNmzl68c8D3BudMVZC/7udZ9eYL4Yb0F+lKe/XbOxQGvF1Dt/T32FBRHLSWUdOB6gjNj
0l6UG+l0kDQOpgA4jmGoaPMPVMI3SPnwLaey39e2ikeA8k5kfk1qwdVpVJvKSqUhg5EkLPOT1xWK
xInx+dyG8EaedlokyERsbpC3SA7+5lZH8zNY9Wdk9Ha2gIeQKiDRgKAEZ1gaJauU9/EESJkNWKwr
H9sFo+iIcfSpsJwi4u/QZb98S4KB/4evUrJkpivHFSIBq+7mJUOth8yRRUC5wzuuK9X10hL0PxAa
lOOzmzI3wor+Xdh9UVUUBqB6kxOUND7NFYYJf7RZGB8Lmv0oleUctI5dHbARBflg+kroNZMPEfOX
RseKJ4ohgzkkSa/daVLL9Bfkgx/LlOXN4uD9rt/uZK5zSXPiJPN0HIpiCTES0CqNMn9vi7d5ipLT
BIf1cK6i81yrwUfD3V7ynf7sgg4nrcZGRieHq3tcCPg8NTHoGMh/qJnk5krQxBvoyXqYObD7TMs3
3LqvdaEgnQzLkL7/WSkKDpebE3S6TPKl/1981sc98st09F05gvkwRIJ776i3h5diGq5KMlYSeEB9
qmYk7Dkmuexuul9nbYYk3Wcoi7JtyghPbJL/vCFY1l1yW9Q6PS6cPa45K1bqw16s65NrZnmeaLT/
mhEHdvJpphT28dW/dZLn0dcwNYtT6wROneYN2Kjpb5hrkhavM5jebiKhsvWVFJpqO3s0Vd431frF
bDcsHb6ambD58wKpWrkSn/H/yBWAo4ZpgV0A9do+2h4UkTpVCFqzzBVitLx+Sbo5PBpYAVkuXwdJ
rAIQv4vC+RQuMrMxtS0DeW7wHUTPeydgQHozMzbe0N4ZfJh/cYao6DEXtt3NoM7BWCtNI3bVJmAh
VsZDwp+DrxY2S6MgdcPhrgSupt0gLOQQ/lQSmxrqp9rjJDECWTqmqR27dh0lV9qsgk77EQbUyoZA
imHFuM7CIfGoxWWQRejfmaSjOJDz1ZerHqayWpH/qCopy3QdTAN8QXhpw7BtcjfPpjYHQM3QeOQ3
ELd9oHSnR6E3r4bSEra939mrXewHYoP/7AJT5BPXJiZ+7AYvl3AixzncxUmY4GvfoyVl1Zt9Dr+T
nnMarXn9FlSjJxmXiyl++2LtVV/gILeYfJvxiyIkTQQr2YzIg5mQd7zpE9HwGXESQ5Cr6EWU9CoM
qkIIvNvw7zXagFWeZlHN2CXUlMW7eptTd3YUREkdfgVqzqqpmGakoGwR0Oa9ZFVshDo5IUbDqcaG
7JsHmc+DAgIfz1v2/6lsFvMfkxRwjVDInji9uUdqyN3oU7GycP9ft9ZbPMzasUZzJiMAJkW9CKdZ
25wJ0mNnzsI9tGCLzrutN5hZKy9mH76lYxaoeQZlKO2QK48ak9cj7+9X6aoeza6svDZOx9D4vPg0
899d4kUb3pH+eDYhYrcNBeYu/ofKuscHmYVBWTl0pSeZByqirqVo2rQFXn1CWSzIy2fk43gQ5BnC
PfdEQFqZU1FUHAJO4STT+92xMjzmz9Ngq2zQwuyDMw2BMV+G8IGwksVXiYWyrhFD9nklkwvw9mpa
rVvGtGZOfYypck6RXtf+Ls5jNNWmZ1TqHTj5ZwRZ/tNtrQTgoLg2ZCLbQlN4D6KnmqsnFM/EicZU
rEtGtwci+zn4g21L8LX1lMlubDqp/tq33Vkwps/yHRO50U6iZXCSdca/WkAI4nIl+A//EPfi2zE1
cxsLF4T0qoogXUjKolRkXxgTFZEK5zRA18ujHVQL+nWCg0U0yuVcm4dFc8y+c2VSutHyv4IoyUsc
KSX75SB37tk6j4QSkXLpQM80XUnnVQK+jDu5C7IfiqNct8g7F6SonQi1lRFSGX/rrzwCyHthjeaf
hS2QOVOpbxnKb4EjTFoc0s4qKv2xx94K6VCCx0vsjaeDkXelW0wfNtJXhpqU5Q7t4QimPSr8NyMt
s3bFk7AH6dwYZNN1fXhdrkGOhD09btLxX7nr8HVqL/eUCZAADPJ/kphvdpIOvTnIn9y001Z08zmK
5BHbuNWlOaGMz7S3mnGkkKfwDdHoTUbMDiX5HLI4u44nEgUQfKpRQqBuKyNXJbZezVsOgHJPXf35
EhPv564715kf4Dn87YTArktpCIlw7KGt+SjyzFOwxqTAXzO9yluxrU5/XFMHucQ1AF9II/7DPdUh
waOxtCOaAkOhEcYme/fiNYwTBGAuaVCCcBsVvxEXr1KsQLBZUU/ohLHmdvjOZx9vg2Ba7DO5XV7D
F9B1BGsFKW0K2NtCPgosjPOb0i0xbp7oIWC67SWIFLHMV8GjdVRDodO7pPIE/PhkEBIaE4FkO1Z4
pzyI03LTr8rAtRdcMML5vf/CF8LObgruco7AcfJE2bPUz+y8Igs6atSTOtZHgjGhKPUJ1Af5dlVF
W92upiL5kMdsjYaxihyUpT8x2zxirckkvDL73hkmNqNxsYeM9qCb1OCVbdmrXAAXB0iYGi3G49eu
BonAJdsrrm072jetPoryoHtlPzHsoaDvYxtki+WkeyocJwGKEAtshLi+xcTZ4bF/Pc34v3UIMr+8
H0r8nXm4048tSospwHokhGinoujjTY5bWj5x4aRGiJIvt49RsOP2y1ZOJKPLwdJP1L6F6MRskaEM
+lf5LO41jKc3/6kSU+3VrvN85Xc4EWx55k7tismWv21WzAaUIS4PHDPfL1ZT8j52AOwn/Z82cP7S
PzhEOqnK7+mNDLwmu86z7i5hXlrF884q9huAzWk53O6LzbhExoyGSQh+zJLgsg2L2jBIGQ8MQM5Z
35pjCZxWgSdCqt8A7JLbVfGf9HQkkWY/UNkcg6e8262lVZU0gRsb5vG3QWw0lQX1FcJGdjxy1gLY
kHxj/5xcHMZ4tTxlzUd5eUGs+q2SJiBe+dEAlh61pPiqQAfvPyZ81t91jTbuvungc1YRTj81kHJF
X5PfnuKdg8cydhY+6Unn8NInKcIaGKCaZWbUEdue08/+e01eofqj/lXqDWSxhss3sCY8z5h9z88D
9Tds8LVZ3D7v17pNN8jwCbMwANlfkBCCqD+FUAK34iOQDJamUkOTEtEyrzGH438ISnCUqcGMKAB+
sYWT9T3gaXwdgYy6aNm5djbf6MrU3KeQLZ/3xqjgcln4hJgud/O98409vU3vEUY5O+gR04a8qQdp
IUwiot2RNLRIyEsmSwTmXtN56FAakBhIqQMOYANO7qjHm0KFYLJ+PVl8nrGR8o+xlth0wfZUZT5j
htrIGSgLFYSm6IXfZBGOR9MSD6NzVSF+7S5CrCCvzT6dA2WLk1DNE0yEn0yq/j2Ee1iNHtbSlZQW
O+c6Mb4OuH7BqfF80sAJuV7+qqjHenWZPTV/e2rBmdGQpEr8Y12TGgwuxJGlqIvFmmAXldTNdLdw
mRjJBu1XIonP7dGVO15T+a/hovw8/GP7m5tMiTwWNWLFzGMwGhnoHESwpAZwFV7nPYnbV/Qo3oCr
uAtWNgemaxdFP3nrM7TvmDR/Q5f8fRLi/DrWId3R2gbLodQrYzAw+cKZKHXbkt8lZsh3Bz//7a3U
r3ylb65aKb2tAQ496J7ine1SgCdCgSeMVf7BNt56GfIlrIE27yBZ6Sw8Wq7mIn1OdrP/Ze7cAEq4
/u5eqiyorrDRP4u6JiIwCdxAQygjLYQnFNl8/fQNVj0lIg0cGqxdL3giLYUPj4BEGTFrRw4TGd5+
hfVSiJ6oiAf6gAcaDYB81LonK0lVdbg2w5ez5qCWxqPeiqgn2tYF6DnIOSI8lHIVjUvcow5oxpft
hHO2mGgQICkqQKgxKamUUi8Wut2pDByIDmqGyKYgbG3zXJNWT4CY4i5tMErw1JUGEO4IWtmmjNfT
xGo46aXSGh3Ik91ttHhDG2HcLgHl9nqP8uutcPA/7MafNJMpGShwoBowFE0L4LPJYIe1vIF85vvS
HAMEbVDMB8BApuovDuAJSP/Qy+N5TdGp8a4hbEdOjm7LWL1FtEsQfFVrzWO56MsqdtGaQAFbVmxO
iV7SBXBzkSWLC181+mLmMOCDVLXUN6nVQWgXfZBn25v346MhCxRARtAmCntmRs2p/YDcFtKNyr38
DXNcPpi/E3bMMnvkASxhVgtdINm6Gx40FVksHEX2tv5RODy5e1Xamdpb0vxq6Cd6Y1+x3LcMBTVg
3jM8NuQdnpvAmdzXlrlmM9DFnR1KUSRVSwX2Lp0iOTy4QO4bK4bZDnMYcEfN7V994zEmz2xMclhi
8hI0JDUNYfOZ9KLH7vKqOnS76mUo0xB5lE0IQDokeVFx8np2wyLXXsIjuRVxXXeVowmdJcaiPxjR
Cig6YZUngfOW8Lt+AgSogfq22h6VCyjL7e5EtpzUXNjVL3i9ylGatT10nIZJAJoc1nXmXUTuwI7h
bhvz7cclIN2NePJdcNjFLz5aPbELZ+HwATPo1Jlg2ySaDEtN23LS95Le5e1XMK8SlzkH+ykFeVJx
r9xpkseIUcbLZILWi8nS5kLL9O0ZsZxutDg6jqYutAa4Abgdy6R6R4rL+HBBQAcWIkdQLnwD3wfm
isyP0/LhRqxKqCIlr2X5tUKrCDUkeMVgrZY6RLMaAoJDAHsi8ZCG1/XwyT/zH2A//aJpMgu9t+yX
oS7s20hOSXB786Rmo0PZQfmPxjBpUKDMbIgMl1KsTDRdfh49SrCsvnvXHkeIJ9AAmac+FClviSxP
QR++a+/5xy+JZVE/pMm17Ni6podI8npx3F1UY5Idf+J87FINfAmizoMWqBeCzXSjFMwnKWwE4XOt
kDvYvd0wxmU0jf91ZEcEPtLKBsg3t0pqEjnOOaDHKMKFHW0XxDC/mf5oBwqm9lXO+2mLdhxHesyI
kWJa+rN1NG34tGYYIf5GVIUT9hDYr+jURI+2Co3NBYXQYuZNNtWNBomE34GhRkJn10RIzgF7iJaD
sKj5lRzA2NAHV/YHIzADUcEnkG9onE9NKeJQkWDss5QEL6j0w5QklB0qSrLszPZ0cBuLNKMwXO/y
Et4//qpf8wJCm40KnjYv6I7oqyOCUOiTlNIlkt61WX4OOGve/mN8kZwpPArfLZaHblVFz0Tk1Sbr
YZJauTMhd91UofGZxSjv0tJzR4dTyKMKD8CAVpCRxmhv+qsKRdAZg+/eqQvz+r3Iltn6aTE79hOO
2aNM/LUeRt5mXv2nVpTaixY2wfuIU31ifMawwetzEXABAyvDAOeg3uAoV1ylMoM6DFE4EPos/akm
SYPSY3f1qIulKM68lFJh6IPm4aBuC9c+FpxNHLjSMlpgXxKlKG4+4Tt/xfWqpTqatf0LchMYolsV
p2mp10PLKVg0u3jq+lDetmMuuyjhZQA4pyg4UxAroUUTuDuovDljrdf9IrMlpM8ysZUbiokj9kjR
DKgxGc0g+Vd6S+WmRcFi+NTUQqRedrL+djxBSMMloDp6Q+whQDYL4sGAdWY4R9PGalXziB6KLA5V
H6qa2WM54tVOP05aRboxN5507L4Kys5kUaRsl0eW5Q4RsGGtulFhLQamJWVC3f/lP1yVnhUYmPeF
xIOFtpHhg9kZDa52pyaeMJF/UiZJdcNLURKLmCiDSYMe7WQ6viebSLrriSRQzQPFWhMhqt327MRl
un9SqOwzl5d6Hh330dCA2rxyu21/LHcKRDfTulp0FYCUnqDwKXG1B8LoVhwVOOARjaOluDpsiI1c
E98YFlhItodgxcVySsm7tX8FG/tTaBbvjak/qnGqtEkb2wCksW93BvHRv5UGFQ+7Nqa1VVupkX/Q
Sqeb+1s2rN4Yc301p/2iUSD4/sRjrZl0Linv6dBVTOeddstsit73g/c7CGeBBt/xcAL5jtGPVk9n
NtqQHoEWZQay0cX3sk5VmIsGHKjZpCMLIxIdEZu1taYKQeOcarr1X+UuR+bHMXDe4dopINErhfyz
0wqo/cIXBNEZgmcAvouyLLETW0dS9fIU1FwlaSuANn7Jw/lQHYuMezPoPJoQ7kRU0JZGfHCtHmij
24AFDoJ2ontvqyG/3TYmvOHzvAKy2c9REzoSEs0sBN7VtH2GcoYTFBJ5YcyEJid0xvhm4p7bHnXx
IAyNF/2AonHyZDx2WKHWiaWcxokkUYwgg5enoYfzLGksYp7ow6IYDcLXvCdqpeGcJnGBx5cR5NBn
pfkjQQ6VFgYKRsx4ZEXK3K0IxHQ+FQPstnbS8MY5j/M8gfQ8Etu53VSRNDIeRDtIQT4qOCKvFAwY
dOwFE5B03kIfKx+5nzzoT9wecJUnLo6J4bOwDSalh0i1iaILOi7vVHXx6jVDYTNut1m0w9II8jHO
sHFttStapApCjnrsOP0mYGmmPSbsbi8UoEokPGc2VpampYf6yRbAesqEHzOpW3Vr/ZRzkchMb1mP
1Ffdlp+FxDKS9JEZWh+VU5LFo7P3jISlHg4oAjiJrSADe+heHNXYOioYL9JiqU+2GRtfz1EOTMhx
1T8uKhF1taWi5a69XZq8VQk4/y4E9yxh7isHgEKlIqrEd4T42DGK/Mx3olIq4JUYdP0rihZA43y5
9FEiD+pIFFLqnbRGl42ezlDn1Gr6cSzl1Ift1z63QHlnDoexN8r4ER3zl8Y5NlPLtHDk/yzyxXyx
Dj/ED5P8vC1q40nJ8niRwUNvz4AWY550r9x4TiJ26RgckFJHRTcEMfqd5jrsJ8Pr0NteliSv+wAI
R7DMaGqjvrslZ4ck77ALzdULnZVfYTalvIyLb3SGZUwvcG7ooMGV4Bw87GDOj3I0aXdzwHe3ldFj
p94QhUS1c148z9o9FDG5GlZ2+SF4+DpFXYkKwKUs6HbYa0335n1AxZazowEaO9P5rIj3bNFAd5QU
JebqcPYQYXs1beQ3aFwcMeeSqDIHaXxndNPmdW58OwqLOze3nHHNiHSAGcpbx1QLEFKt2isWYefP
8F8QMtUs7i3uWkyQ/AROmrLN3hmD3LB/xD7E0uHt+DfBFHhKP7IWgJKp3/VNIt5sxKNQhhygxE9h
7w24EjgyDUTITmNuVNXkepQVA/vbxC9twXKMu+0KwotALCtLeBIQpAWgDv1KvF0dZLYq1Bemt4ZE
RgZOuTmuCoMbD0S8XzexWVpyHeT3fj9wmwHo1Sj+jTVJ7hk9k/LISfb8mwgWoAZ2kqzsaYxsZnqb
ZNuRT0yUJ10mcmtCNEd+5c72cx5FShFK67rXYmkUEXmIBEVbhoO01MQjteWwzcicWBl/PUjdjwgt
p2PiMX0RPixJn9NoyeQDKSNAvP53LC/gp3hyO7TskiwhW7q6kmSLQBu3fA7wqH+BCohh+eC5OUou
Jw3A8aLkBs5F4ydYeui9fOfjzOERI6pUQlkG1MJtHcnPnw6FiBxlNxTdi5dqtuHg5QRuVgbi1L0D
FQR1l1SLclws3MeLK1y2W1lZDmH4aOPA9Qnc9SQO8u3VqnfGj9eO6bTD54Zc2immyRrve8HxUZdC
xjxbcSMysi29hWvCRoq1dRE3zEgwFsLu5PCELAZxMZnpmKNNKtT1adwORVclqINO5cn8sz2Fl4sS
IuLhQkJkLWwxKztRvVFH9h5VTg1gQrXOGp83kJJKhl4ZZI0bLVvhszZ1OLO7IP1QUc5o2ilV/yJH
xRQcP0V4WEQx874ChlQ9b79/1WpV+MlM3WXeqEBmTi69TMDc7RFDlK6zrzglwHNhQUQlvw8BBPD9
jAjDQPdGhB/WR+wov+waCdBBae5cW7c6Xg5TtEtnSw7b3cOGUPTxTkh2HJiCjGqQCVNUO8YdG6pC
DR5WqULzE3hGgtgxP8/WTbxYOXdAorVReEQ8LNCsTFJMiBC/L4QQLPSmJcnVg0Tg4t3c2JfJhJrs
WjGKKE9VvGeghR9YGbcOPdyBEiojujz4S37KjoQQKpjHlGE/+y+WQw3sCQktpccX5yfD5oSwm9yi
bPtMO34q0mwBceEa0RmR3OiJXIbOX8aCmPH2GsXeIBfMxNmEDNndi7+P3K4WqQIZAbFMfCZ7dFQT
rmbATjJ6YUesMBwlAR8b8ULmreCYbNLgZgI5mHjEHOLTdx7bsf/GlrXOpoWe3/z6Ouib8Jxw50NJ
kJQYnUL7mdDaCTyFiWEEpLg2Lsa9liF3jti1MY5ratfW/TRD/PESlmCpcB9AfMotCgyez/rP8CEc
IkbgCNRXewHlOCgPRQc/g+TulHVyEWgQwEriArNuH4xbX0Hq/UaswJ818XVE9dmWINOpG0Ut2mp9
Sn/gW/z9PEVRk8jqT4pctC5iGmLqP0CfAYsgv250ijZvLHR44gLSHCMtyuexkH9pYMXAzdwdc/nt
BC1GeKKk2JKE3w9RzNe8BxEPYyoUc/KzrzlKtUfa97qTe53x6/AaldsY4TDD0l39e8UZ27hB8lEc
IMXwkDDRKqVh4mwxGtnIYQbKKQqiKw24//dU7xC8jjuaJlZ4ZR4B90y2HDH8+DdEBwVXrMdH3qO2
HQMongmBf2wUY+GPNlod3Sfbt4sjo4vOeZBYV2OjddDRk60qMy3WLaNHdldI3XreaqtXyz5V4dp8
sjs/0vBT/ruHeIxkb8wAGUZoZuVUSPSS6IvLes0KlYJSFiXWxKphYHBrcjswcKaDc19dz+7kD+pS
JgAgN2PjT/B4MwXpm7SepdNbPkGCYJzW3kbJM0EKoVjTvLXhzAMHm2i5UYc9ZHJfJJX537DFlMHA
lr+44/QVPS5QsyHwYhBgENvkX/QoiVPJ6Aht54rXpu7WqmI4LBG4171wDChWJGM0ZXCcwYbRvYRG
gCNKVdjV4J5PxaCoS3MCJ1JUPiaLd9BWqCPkq9jQtWzA47zpoPD0DJrNDZINQZ2pbNEfDqH2VZ7y
GuxH6ZIbvDzdVJWk+29n9Nh3KzXj+ZXTdTK6O/7PUc1eL3sAlG35E+A4GydzTnukRNXUbUy0HFZX
LGBRitzFtfQEaC2jZyiJC9HQJbopDaahNkIAKomY85Ky5a89a9a1ALsJ+G7zRfSaPeDQ9Qtw+9+A
gJyQ8Fjmg6+JFGMBT5mo38rwFKv96ITgrK4yAbgu6/MfYuGSi/2ir/Gy74qxDnJhBPvRy/teMtfO
G6yaib5DV9bIFRvgk39Fxx+93fXPy4LNngBv1ArHmY+PmFNiq6Yu2FSxnTmFjVaFRBT0Pivtsyis
TMm6HQMZWVKn31kbVAtUxAakUacnaCK8KQHUEtC5yGgPudQyyIoZTv7WCbhTFNzvvMNuyTKibi1U
nHPts5PcwA46Ws0NOq3EcY+tu7TIIsgkkag+UYXjLDIVwjGAsMqdgnsgTH89CdSeKeN5z957LxDD
fy2qSg3JB6fYJTL8cSBQq8YW/cWKEPgaeAdKAl7tyaIZd7ZYAivXR3kRFF0hfV50pxeBUoV6cco3
gcQZUSTVLdWvI1H3pHShFOUVhdb4LYhxMbdLFk5taqvwY/Nh7gygWll8wiCKIu/+qjFXomQn5HAS
8H1F4SZzEW9gYkQyt/0O6OouuB8WPgW7tvQSRKqHPCmR51M3PIl6UOmEiqX332UOSG012gEs/NhB
osyOLswpTGjc+fRZaJoxSR0s97QEtMz/w6rDehxvXCvHRR0ugFW8wHBVjA0SxWPTb67wQVMwnQZ4
JeEXpp0WRcGdyYtysrHt9OoLdTr7IH1I26z+4qt4YPceWDrQosWZ8fkRICl70ZAidhY59qHyUf+C
7wcywMhdE+yPXPCswI+JI0Pjfk1sHbr5U2hJkqfX7ABtv+Ss9iIx657jFd39aeWCCKvxxHTaQBIq
MgVMEk3w6FbkkcDaA2owjnkVdVclFiftaYYH6FSkHf03P0yeM3HHnmHcw3MF7vAON30GjBaIktCM
tS3PQuJDsun/LfTJ9tfoZRAkm0gbacuSHtbg9LZMAsJ+odKH7pv3icBdb6oA+FkzgdFC1xLoNrbq
XhDC4IwAfAtByBmLqFTgec7zoeqpTgQQofrTOJ3TXFSGTFm5TiUIKmBbxxIrHe+w+MtTt6AWygj1
RlaN71eb3fHcj3KF81FtzeZjiA7tBTgJJMHmktucQRxssTYuwbO8UcdZUfm3celdnHi8MxOoOyuZ
OPKWaJxeJz6pshvCDr/cfep7McGcvKyWxsGqJb04Ww8WNLBG2JdbmIHDP1wqxrM01aBUPVNtOedi
csrTPpZpABtHHwgRRpOQUXacwNM5RH8ZbwuEsKLitHPrJPacbfgWOmf3g6PIRnisBerjKQMvIuZl
9umR9KdxRdUDGLt4wfjBIDp/crBuVDq+zDlkK77TOCgTMTXzToAeXN7f5yoUAKZ2Pp/iPPLNKfv6
NPU+NSI5EKFK1oj732qiB3AeiV/MshE1XT5zpcOeTFAaozsSgt0FjwgoJ+FQR/Jhz0KwIxkZCN6x
+tH9Wd7w5vvGK6qiqh76QXYt6WhLAcEhGkKkvoc1h/oia7P4Rbpmqu8YFw++40ayrJgQ1gBkWcUE
PY62aCDmkYav6gREQ6/C8gDo0Y1FGJXhMVttp9/LJVrHf5M9+HGUwB+6bh2E6hEbZxcPUB2chK6J
BfPKK7o7P1mRWRcL+bxsdTwDwB1PQ+RzN1icTKSEMSAKAEtNRFA/amDbwDEWDQhsHhYHGUrL3FvO
HBEut8+9fM67UiKVf3ZEZ+A/ycu0vReX45T/IUGYpETM7jceBp3dV4alehGN4OrrS+QBaZYPnW8f
Rw/Oi+MW50eS/puSE1wslgxDH5Q5m8+41IDsaEihm4lcw13Npd7LLi5Im0MrvTPCsJnt59pOockG
lz3gbKRH1g39VEaFlHiKn8laFLaY+keoa5ELJTfF+RKwHEOEweXsvS/eI2zqbzUTCx4HOdbA+y/X
N0xYb32bGa95+oLfjckjGyEIRgUv4suCxaw45cHrm755mzK9cj17ymIzMKODWjI7i/SAN1+x6zVS
E8qxWd+RYLaTi4anFM8crgXUUfuwtT2FbPpn1fBd1hzBmFZuaSh/MNewJFBnFBXVt/RscOg1AoC3
dbgHZ6W3k3J+94DkVcYygZI/9gEzldH8xFqw44L95TDAB7cYlYc0e+1ioxpD+xFx/5XxgXjwiWfS
m34tE8Ke5CxG0dSTNNY90EjmoQpWZgYPLpch5o1vTtwSRtYkPIKlJ5vRQ7faeBYQO5pHGWLfV85B
weo2ut/ZSwYgJ3T8He2PuoJ+8V7cvnYInhGD/CCOEwu6cyEluq25u1/AWEsGBEPuhTKHNEL7BDuE
5gKNDSfdJqfVQdk79MOmppW7spF7SXT/6KjscGqIO2FV5+mkvFdZyMtUo3l6LXvAwOI0GbX48GL4
f/b49Edg6+ZNE+FYnyHhRhlCArIlHlO1o/Zd5vYAPrzOD107n9foMLWOhNBBwH6ntNWcBNYMWfr2
mPclnAGe4LvLdEFOh+1nD5YPDrGhHxUxulMAnG35kV5fS+TkvcicNXz6awwUX7ZmxVE4p1XbERjh
o+sWWj6/rGKSoH69J3cD1NCB0UKGtsXioeOQVtTk72LxcQbwHW5UcBLrBN7zZ+IvVj1lWCFUEcjv
O5nbjCQutKOKw9GSrMyFBoY4Fk9RZb4c5wJgtBMwtL9OybLciyzu+q/0K8U0W4PyC+rPq/2zJyN4
jb06wPIZIxsN2DcztU45zjjBEj4k30vZQTyrIQtQcgAgfXpo7oGGoWabSo1CgQ9ubYBlJbM1jvTs
0Q/R1fPBuR/9V7qOs9vzmN4vt6/1bt6mQx0UiyI+Cane7fD+Ui4KXSsojpimmUV6T4nb5NlD+pXJ
LY/tSJb8r1CJCWXE711bjmSml++UGzFtPabkCUxL77lpMcV5BaUTKCzBMmklsj64MZHJ8vys6px9
uBFCTr7KO3EJvCUcyXSca8KcDEDGEv3iSBOAl3M3V/nCQvuE+SqA8KbjSP6wfPnsMYI+DK32Ase+
PErFBu5tgdN7/QsAv/J6/Lg7pkJHLW+hX6UsE5J3YryvxhF5eJIrspgFFiclRXCzORKhDXmO3Z6T
0dZxoHwGFiQG6iyy4M51SXQw9iiIInA59uN8VI+GDvdbwDINHfW6XD4HfNlrUL7GuCMsil1qbvqT
A+UbEEr/Iz9/bX9Hk6KUNBpldGbjF7WVkfUaUwx3jiSP9bAQmOY6l2tNIaiHNxSkcw8Pqje/wADW
6byCq9M+n3lI5ASgrYsdQx1eFIRtBCo53rZjWIm9JxIdBhSBs4EgO9Ud2GjjQVzcHnO34aUBXAN5
iVFtH3Dv9OoKih/f6YzSSE36YU++QrGHfuqnJz9Y9mDSiBTuIcqVCqxAHc3Q8Ey/Ukn286tttpsG
uhzd/rOKef3oVttBQxxypsp7un21r4GY82+RkSQah9U5sx51mPe/fd9ZIY5ZaEQxNW1A01ph4yjA
6t9r9PhLCjxUX0+dFVjRPOudDJ/uDH/9qiM+ThnvAjRM4pM3ympzgrhtOEgTFQPjFxT3vr5w4AWu
eQbswp3mL1cJ5eKVJUFVi/TDAeRuB8IlK3qKoJNPDlOTjeytF8iB9mtCp3p4PTr8PZUviNCKGlXh
nlZnrX5uzrMgZQVr68fIDG3KLh6wS8g4cuBwZWe5Puy4ml8Wm8nnK0rlF0aSjqXYPwlT75b/FHyH
v/zddzY90MxcLqjcnoo7MVOsbutakWZ9IyOmPOfdUBFWL95H78g3WT3PceTOY0SlcK00XCgx2aiP
dgeyr/tMR11wpriEOiFdyXCprSJFzOsmpOXL89LqRGKLs8vt5WMaIzTUrQnEVOVdAnhIBUDmCJGI
I/K3CBvR0PbNUmYWFnMe0hzueoXiI7cHI5XJaxeKgLsaWc/6G/w8Pt2yoSHHLXVv4TlcJY0D4Zn+
0z+YELY341VPuyZoLxGjzHvZrgottln2qpJ213su+BYgNlptzYK4/cB0nupYU+skw6uhTHO/reG7
w+FbdY5dXmP6/bImcIte8J3LIg7KB71/662rwtncCy8DQ0P7FBH5gLSUqrFePHIsYMQ6qz/fdFWs
qa0COK5sSCkSVeD3vaB+YROpH2yUDiTkwvDPWUVBAnYb4bYMsJgs/rNfBDLiixmNFxxolHetY5C5
jsl73o+UhLiY/M4dZOOkBLjupjm3JZtVoz7cE+oUAaLdilIWmynWKnSVxjysuGLbFV28f9UD+3la
LZ9WlBGIFlkIwgpbPYkpyxDaKc/BaQTwWVU60h2P9hKyoDNBEr5047rdh6lJgvsl7S3zjZZ6V+om
hyXbZaj6Cgi/97OfIa5yHGbLbTZZ4AhjVOWrbWK+Bf8VLSyv8wKXGPZm7/vTRpxrTaMCjorzzAOI
RYuj7HB6osrZJkNmY4Z2LCXl5KoxoiLMT4PZyyxRgRu+iCrMajAYtwc2767f3uQ5yl1taLuj5caH
cKs2x1UhhSswByzvPtwkdILYUwlOuKejKTYZPErZAIVkymWOl0bAs/sPq13KubbQq3RvUD/y/1na
g6mozhEVC7HNIdNH+zLOb7N8AWJBjMTd/r6VMbWZVkKskh6RAUBptINLoAQCMgCLztVBEJQqDiGc
StfT+OsCD/R2OeFLzt+m3UZVdrED3yoA4KhvUftBUKZHzLKNtTC4oIAZi4TN8Vu78uyvvxMj/uuk
WfGslA+5D8BCdAmtXghE1yBkQ4P9BkMBQrG7xYa5lG6YX2scCChp4wgBipiGMnkMDYGMSkGWjF7m
jb341/YtnouQfdrNBReSR9lRQlzY62biBxT/YsgZp0F+1BOdIdWvI0mMj/G+5fCAdCMKN+qg+Wwc
YmpDbwb42VvGSFgEAlZ4/9WlQ6g4neHOv9P1wpgGWuI5IZ/H2lNLbkS30o2caaoOyu80CzEtAbyQ
X74pVk3HjOXZ5QQrWg/vYyQuJ9Vf3DVv8BqFchOBZ1yPP737/zgvo3vRP7caE9gVrWyTTkGw7EiN
TNaEzWPWKsD9IvDWfzJ8loFgLGrgOdmI+CSjtIR6jg8dY1ddUR1kqPVlJHTBgzXu67x9WeFusE9O
Ppre4fwqx9KWUpdFIqrIlVstYvOrgj8XlpE7jhO1fxN4VZQvlDlwYYRMFKf8VmQOqXSoGSDl63bf
YhLecgxKOkxAvZ/96fs0KYF1qOwNmUpI8RN4NOahs7lMv7Eg1oY9YMuE8FXHv2VeCs5LTrQgBEBq
7YxtnH158AOpY+krOPRIli9xSFxQjOuWNhytMdTeEOHSTX7h/qCllIImdofO/q7wYy/k066tusTi
TzV0ycCClFbfK9VGmyFxcXviWM0+zX9WjnttYr14WpdzQbr7ZcetBj6LUhN7v3/eXFJ0JeOCf0Wi
xg/1GJ+fIQVVdsWwkJVFG+17n+cw69M4An+BeSxWVk7+PtJdWKCJe21Jjg/YioWNto86unV8WwHP
OspsF6ylprPQxxXMTBS2nfRAevOAP6xiQLVD+ZTXnooHWnNO3fiKiy7sInTcZpxh9hd1A9ifsKJa
I7QwqWdjIIjY7Qj0hOYHG8FM4ZKN9CfL4tdRmo6wLUL+SaII0FjpeHqQMuTljl+9gudsDRL3WkXo
hjmH8vknd6bqqZbE3VF98PU/ypn8N8PfjCOYwde14F/PEnDzR3p6w5Vtv/YG4ZJ5TqQ017X9+An4
UhY9RmkfIjbXZ41Zga4MfWw6jN58oSoLGlAp00GqXhN9zgm0+md6RXxquoq/jHqvqmV+7iNkNbhz
QhzPrasR+D/+Bu5zRYvLZuedCjqTDOGAufrRhNVufB+WNuSvZHzyM60CHEVRA5oOXopMFpKxg9BS
JlXYIOOEb3YIpasXESqwTjbA71hU/Bg3p/y2BDAYh4ttlPpS82CHH98GycxipLZn3fn4IXrlhpQp
4Ned3Uo0ptuFryVU2Zq4/pdIk+qHp6lkJQ8WkkYSui3570FdD3UuwB4LAN4aIpDblSnWTyHhFFdo
8f2GCtGUWYKfq57i2TdkKn5z0jTilWYjGMGyxBWVxhSux6TcXY8N0hjrOkUAZNd764rfubFawikK
OhVOrkgjaI4JUqLjIuAzaLumKlHASiIY4BBJrXSz4/9zdlKonz/9BNbDWRmKA92jCiE8lxRVoVIt
kqygY8z5l1n5apNbT4RLNhEiF5ohpYp86R+RUkoyGv0BQ8G/BiewULI6sLlcGzALINlu/rz3ytwp
vmrA7St3CPMq1Juxj31/VcsBgoyReokCNKuyEY3Xd+3drE3lgXtphfRH/pKMkUB4a47IAEDoQDck
83EvEKwnpZ4BxtVNN+pR9+K5E1PHFl54S7LIygx96ITcondbsQ4EHvV0K2d2b+6Vb7yoL70zTBxz
KGBS/imdK/L35Ustz4ROlYntk5d4I7u4Wfiulto8GxQ2QCqFRhbzgIFLO2FAHWKaaVU7LPiaXmOU
6wy13EvT702nqHoNGuTWklkaXVbNG8AEgeCnHL3UH1P1XCNgQFWnnWP6d734rXR1trbxxHgb4ERW
Qc6yFrC/+i8lNYm/5T1fWmXvs29VRRdgb+/CSfzkygz2aXpDRCtrOkUw7GEjitVjPJFd3Nz+BdwM
LbBE1LKwCGq1gMKOM9nj7R6zWwAvBB0c4J44E+7Mubv6c0U0v0r/adROieCRp6Bcn/8tVqjkGHm8
3zP7YNKB6tUt7+CDHuhmVT8FF98OfY0+YVeVz8ptKMSO8MMV8iSbi4XbLz8VXAQ1SqTb5W18OvHv
o8r9W5IzTMUfD9x+ZEOviXiW3m4buw4HSVK+Miyjt78ruf0lNE+dnJOYbonQYUVH1oFbXTfuFiG5
zJrAU4s7VDYPfedearXElHxJq9F4lNZ+0BHH9K7/fR64SlxXaP2mP4s4JGy+IIJzCEOrvvtEgMc5
oYt+SCC+cf2BXO3SM+TMepvcRbOtkOKh7Aaq2wN38oWVm/QprajKOiKmxGv+4dNGLOyKyOzyA2TR
5qitdxwfpETREyiT03yh/bfqrxdGWJaf534CUtD2HNT/hrRDm8XGTzbJk9Z87chuqaiQsMNVVmZb
dxiJl20kKhqG8p2gIgjhVUB4lVNJz6KqDFjZVkjPO0mqUezHrrNS7fmcG5Ne9cH1tmY9d2PFjtW1
BUQQLtoY1bUCHfzhM5z578BfBGFz8XKcmtxK3B7h5Ic/G3UfmAQIcionSgZ3U4zLXqvgA+vzLfKu
vVi8PQEzBaDy8PCRb3xcd5spiltHQhQykhl9SGnhU4DsK6O7mQbMXL2eJQqZD5rD3x1mDr0cv5ul
udkUVXFzJsW3LLKhL7uZOtrxmXjA+w5zLQI3WMONRGU40kwOj5uQU8dBlDA57Cbv4sDw8XEcVMvA
pdjLxoyvya+F8krYRQYh4ZeY0CyN9HDeFVFfli9YRI2TwnXmXxCLZbRTgss1Mwvk32HlwButrncR
W3dr6pKrvAD0jjUN4zo2VLzbMtIoFCA7dFMV7GrwZqtBvkAmvuR9j5b0trZJQEyEdPc0dfL9ED2Y
j2aSQVQdJv35COd+8S9ymz76XEVkym4O7tbxFlxsOS3wFnJeszRe+dUe65KzWNz+WCZaZ/cyxyeG
JXRQ6U9yIt3Nxw9sDyYdAJnNMQYfKzVQOZAbiLI4u1yC/VEHZouXdVtqDzMDcUi2NyhOtIeqLHRC
XBqhXfw8YcAE7kw81TagjSnwrvJ0+f8oyjojq5YyYpSkZTQe1wRaV0rbn8iOavXwSl3yxEtYy7BL
C49fLLUSi/H+84S9LV6mF83JCZ8RYiAKbAZWAClO24Yv7kIXJhOXV3zzDKblScq18CNLBs2LAnTD
K1r7VcmQtkpgzAzfTM4Zsy+v98Ajj6X1Is7HEDoM36Bb3QDVEAUs3P+mq32Q0GDxCdtpx1KEKZ+U
rOOYpDeF2cgd64S4kds17jN08688mdVUH31Xih5t/zxhoQXjjqMJTxRbz7xJvUMhh0LojDfLRHta
OyadVDQ6yi/5eM0wBIU8bC33fsz7emDUr2uE3TPHkur5zJJP1cilXu5qqpWCsby3Gh01mrqQi0JQ
uJ4Yxy4j19kMJfXmlDd9qVPxgHOh8oWyDwUW5Cs25O5gyQMpcRtZ/dL8HwQzBrvRlsHQvYPR8O+u
Fzt/QNT+xmozEdesFSHASAvQDo5ejXk5rppQpm00ksuKakzDA1LMhu5x1zaL3SukuVjJXgs+Ad5U
s0Ru+KBcuT/SeaS2dHn+OJXmOK3zJPms9IE+2UwZcRxl3+vYq6BrDKrHJEIXPZAwsAw7Qa+X+fHd
T0iLsYWrlUvQy6sS6BoGyN1VgyEBw3P8qYT0r1iWKIgb2jnhZql9Z36nexAY0IE62CPNFhAUzMFO
fEvULUfxCbUwPh4nhZUgx9tZZTpp6P9m7z6cr0i98ReIR0cwuUaj90YhCcgzTdrv3ugrfTMCmn/7
Lz5UWzjQAq+kNVpJzlLgpM/X6MOJfa5LxZGupvVEdlP/x2QkCrG4CjXwlv45vxzcuJMtFISAL7iK
CxVvYJ7PIXGovGi/EEssAdFCAdyBJ2nhub2W3nrBoTdwcYAQp73SH/Q2gicw8usi4eQKq5H9zQgP
PGphEplvM0KSaN+JeCFGN0SbChrUqG84y6uuEBStTrLjxBqbUhA969FYwSBj4k3bjnqJlvw1NXNB
ku2ksg+EuIfFi5jL1t4+Fi0XhtiIwmTsIToOsx2RMVaEolWhIlsZ4aAgqWCSXuQWayx/kfWHW3cF
1HyhWPaApskWItJd2qdRoWjXa7Ou5GfPxIjXzhcGLsCNbv9hShy7yLtru/yS8ymWVhqDVeRrJ1jB
Ud5QXrC+9wCpaPrF7qLLSSnmOE7m62MdDFHWjBvg900EwD269AxxrcGLy5hv7BxLMBpH/pmdLE4W
WGwnwxCk3oC+4Pc55yzTRfYlXs/WR2UERctmJpwipknPsVE67MVV12czEfum9DGg0VRw0uzJWB5w
unJcbOwpzH0l6gqENxTfSMQGx/qG/WUGqtmDUH9W4VLbmSpOUQIzJyOzJ051J6fr0iL8DivKuo8l
O5IEcsxZq/c+grAlTL5Zi8b5wuGswRhZKI9f/3xjTRPUE/JWy5gETWT1welSzpMM6B0IzollNsmv
sGemrt3659G6iqCbKfB8bmFNysUYyq9jM0nhJKI3fUdAL8rzK1m2m4u5uksUTFK4TONh/Pt1q1dW
QlLxhyPkU/9g6QMtmu/pQwGb0mpWnwW5gNgmMycebS1J0gXWaa6y4+a1BNCyJbqdbHsawtgQ/UuL
N7zLTlSj/wTBLiE4A5385r34EpvfI6nXpfjJBLaad/Gmiw4evC6lIi2hWi7WOLSobviOZ2xbA2eD
KhH1XbfOAh0K5mT/QB49umbQjnC+ql/8mE0NxFL2pKCBc7jzxLv1FdJ4zEPMKOBy5xdWxqOaRbyk
VZRkRonHi2fX0JmbPQF2j0Co7NkTGTI0/519mScssYo94viiP5cz/hHKuhUrDsiiBgHFTmJPa9Yd
ciaQv8gn0N1LGmKP5FpSYtr/56LBKKXOrY9Uab0/V43BvN4K2xSzgwEGEVFnO4qSTjReM3R9OaIt
hoPXNVEs35RIMlI5mQq5EexJPd0s84KJeFrdy93ANVDZcUwdbFnEfXgj7TsiuI548r040AdR7cnT
6quAkjYdBx4BHI0qlvLYmm5EOjL2rhN35T1uef9q5rf1Oiev0aEUcOSocZpPkFs0xDXNVZp9H2+/
6KKZHtJCvK7LLMGHvTbfY3wYlGNTdSZS3Wzbdc532ycj/Uvgw5pikhK0TEPp7UNaQsiUg5tDbxkr
12PxUkkeYvPr9ETZwXwQUX4RoYxfD2DasCdlMTwI8Y5zFaXR9i1FHemIAtl0VfkYBLxqCsjrzwO8
e9SeGHnnxxkTH4TXngBgv88ug19Agc9Ijxg+X0f8cyN3tOiWDdF1tIxwoJ5RnJ3I5a5stHlw6EWu
Xk25MTIssMI61XFptk1Zss8sa/J+EYkt6NybpAMqeF/Kr3lVrXOSI6bNFGHoKwNg+NhO18utbNS3
s0vp13LbR6VEwuTY3mmEo9DsNu2tusxf1PlWuG29gLmeN7lwbBD4QswOIhcP8Flf4a8Tq8b3aGdL
O4PcTJ3u5o7QCfNGaYtM36lNMRebSzw4o1QcqGgz2geoOc/uSMKG5uLM+M873PJvU3Rk95Dkg9qG
ClNO35vJnnBgsVCrMn1ab0RPx0fQuqRooqLwBdLFPIQmus0rshtK4ai4UVaAwX0YLYhfUzVM8/5M
liPOd3+41aUjmtBA2y376zC77Lwe2Rrbw91U+qr+uafMzHVayFEoOMid/gQo/SqGMBUy/4Eamnoo
RRqENFiBx9ntDYF+XjXqUj0IBEIm4N7V4HFGjw0W8TQzQR6Hn4MJChU7g2Uq0nNYWk0WUlFKqX6x
xNUj6k03B58XD2jkiegPU2a8/SI6yTt5z3DWs1xUcVxt2+P1xCcUFxVL8mqva2lHC2souZUT+wvt
2jXd4uqJDJ50yFcfc+cu2YnfSQRiudjYXjsdWel/u2kPUXDuXo5aCKlKGqr1lWK/pmM0mLFIDMu0
1T6AEX456EJMfOIVxGvvzIlB+kdh5+yF0bR+6N1LvyI+rytaTyWIFnEANcyVvrPXFfARvcRIWp0w
qwGaQRSfsA4PNC2VRDB76+LfGe4tNVJzvkhjt0IR1gO1UTlx10R8JrWpSPRFqDE2lQJzXAEYjdrO
ipNK0RIgixUl5ntyA7jSVVOulJpQatrPWmqpzeMKX7TwiuqCri3O3bpQVkAz0XLDGCUxYewmp7UA
XeODh54n5aLpJF5fZyKocy0e005HmtgUrF+7gFrTSsG8/IyzRSrw2z1VLpRSgJD9u5o35X+7zN+2
pihthdCezgF7/KrbCxmDdFvTaKekovs0Mi9tt0ZA5ziP3JckbNejuLUMKreNkH0IKrv6D/jujJPG
6jxoMKam59VqlzH12bnhoc1uWl8JeJJMH6N6IUtOxTbbMocm0UZIcfKoWofZRIcMsJ1/f9Ou4lIb
6d/2n/SIDYwr4Ma/oiPpNvvk455OgQiaX9APt82nYWgWA6PqmpzFpfKv6ylD552kRQS9rIz8SFKg
VCt4H9CWYJbPfZPKhbotc68Y8A+JM3NOsfR201FomeCIAv6+gG7+idJJvP+YQSomdAtyERLnGsBM
by0Pzmf7FA3A9Cgs71OJQ9Ci+/Zsh0y6mgKFn6JHSHNMuivlsucqgjlKZqmjjR1OdFqxdVVis5u+
O4mv3yJnta/X/ChWlmJ3gcyl+AYEQ0qLNKsVE7LwFvSNmj4uThWtVPRlroymrpbq3HW9RCE1cozn
L0okx92zl9mmri7aaxGfcSdYO1jHlsOy4KxuG+f2pFhk96xnqKr4REgPyglogGeGOEHP/UICJfBy
eAbsRb1AK6t3Qlky4swCwCumAifn3lidULfraZS0z+P53g4HiqqTNbk662vo5Uw+tLmKz64Rj+P7
QmtC8Xd2+uVQbn+ZUIFVENQ9BcCrmRvGFDegU9Xxy5dRMw/Cn0jZb9ConrmxbJ+obXoxcUIlP4G8
l7SyXIWfOgIW9odfWlmiR4Qqz/iMPMCJVT/bLi2ZAUUd9/UG6sOyX5uV74stuG+27k2abMtIQISi
6GWxbCmd9oM9QASYe74rFI+zPSro+w6edgK4cIybpn3G5+DAoBorcUSSToHpbBN/jTdugInfAW/o
GSQ2F0i9w2XKOTdBgRk+XhkL0SL61qdoh8xqtWQhuQ/5/Nz1DWY+EneBGg/NnIdleLzAEJHx3z8w
ooMYU4rDx/KKJO3u0DLpiT+O253SAvPgDiIP8zQWQp/5EbLHzNYpmIsZ0B/+V+fujTpIgIDJVf1D
4b/JptTpYdcOrVgpZLIbexJzdUnvyS3/06XuTBx3YE5L7pKEFvIYGQ+cs0u8L0IwHuwbx0GiSgNB
fhGofUUNX33kx9pKOcKWHm7jTYyBemh8vuWxlxjmpIzHisiRVsGu9GCokumiEZARAPgvyBZZpmTD
/cTnSH7EOadAxIa9TnnBIGJXVYWbiUCZGhKZdg/FO1iFUT4G3V2EnuEwysHY/pWfMTYnlKDcX0fh
nhU99hW4/TUYaPvrbl9jDgeSHfWimgY4TLc4ZHY5vluK3hIkrciTgesy5eDR8uCWQRyI+6uCavZP
TYj/Dt6VAUy0HJ7dAliWSfwCTrj8V28wUMqZtaPDtfQIx2k5KIBADrMORS+TNsj8Fi6DnmmLuZXm
IbzC4G7TbL4Z52S1gv0W1lyrkVydUcFerRpIcswq/d7hIEJB9OONTOmuJBOKC2BIfnJtHflMDO7Y
hn0r0gLeIJX1rOWIqVE8kESrSNz82EysZ6wZikj/cLkfQtTxsfuL1toEbsHjLjHB7l7xWQd8+aCd
j15trKkVbMm9MbOCwWU0+pYZktEeIMj2qRL1CniYuZw3Hwiq/Cwy2UOrKDNX2b9aDD2oRA7R3qVw
OQlhpPAbkdTnZ2CFN2dJAObrKjmvKws8RPpqQ9ZmgRrf9uJN0w5TlTCwD07H/zHf6Vx0U8OJTpc9
efewTrXsAEl0GnrhYWG3u/hn8G3P1Ydc9gCjpPkLSuuGsHLIfaF+GcVv9QNzHpzYazebxRLoegqA
D4NW6aMsJc1QdmiCQ7sRpSw6gP9xtbmLgtP5bLsEWJ0Wlx664a1F8d7d1JWAbbgKl+CHnjdkVm0s
hgeauSkpKfEFSV0GgLdsWvP9Rqh4xC0E2carNQ8r+6IplVz54gFzMuGWWvASCXeRn2+SYJ3FpfB1
0uRxCcrTqepuk7eHQFDf6ANh60RwXNudF+L0Bkn4SsezAjdTrv7+at/xUDvkRwT3eoYVFlaNPnXP
7Z+x9aAMUsY3nLTvftV1dOWTnbr+csantn9Tj9VQpChgIPIpfyg5UiaCIQxhpU9r0k54OIXP6u12
z1MK6jyexj8MNeADi+dWW1Ne2mdMN4kwfdO0zsyKsp1F/fZQEgYZehu01nZxW2MojYi9GabDb0jO
KAt99FQgXxP7MlRL+CMV2fkPItLibiTWHaAMvhJiw8aagVhQbFjYXb+iGDaFYEpj3Sjd0nl+CxLj
hvHNPQ9KJ5FbTNbthBM1c/PK3mlqtjqWAlIYudzdHodZmvEUJr9PRx4oHPPBoglNgdn072LgMYDD
oi+EAIJSZOib2799ZGSbuced/d3Q0BgCKKrnZTcC9XIPopNGH2/Kbi80hRfRL3L13PwHER9B74jN
Y5SyBLBcMoLCvSimx4AodOywNasEHTHB5D1B7R8W3CP4z3UQMJ2CUSw5KydP8iONYjDuuXiuJJUV
4CqSz6M9TyDt+4+TIBAVDZ5Pq9fQ8m1NiODbgvAVCfcEoviD+Q3PLBheHQhTO1a9yj7Bdl+nn585
HUdKi31Wf0hLDSYcnPzU9/Lx4rAWBKPFWTalKj+QQ6pCpFVb+jcr6itvX8SPh8en9sEOAc4ewe8X
JxM26Lz0e3EdcW2kKL+gqgxdRZ68Wwkv6KdbmdmpPglMbRYwsDdHCRW7WPNb+t3mjLv/rpH7xGLF
23jxHPfbMLW8TI/UMJaB50f46Pk29rhtflA6bGqi0tprl0YlLgWNE5kG9ict2ujL3x6W9RjbRoUb
1jTcmNkoCCnokye54yoBr+04qt5diFGTEg10fYwXmnt8S++9C7gga/JH+TagXAmqkvE4bevSU4hO
8iPjgrD7iExcJgtY3kL2KPBwktK3GVjDzxu+RqRSQMfJTHQjMQrJns1kY8L8IDZf+tT8u4MgomlR
MdFA3tAQSTArPNpCMMwnVd9XxPTx4W96AMIYQ4jDo4CeDMx+HzRgEmDX4eI/OIYZazWo36bsQeDj
9IZRdYW8+6eNk0ejAxNP3TzkUpiZWZ21tq2CP19i+4eGj3QTAbJEumTHJF0WXzToioC5J1xJI84Q
SwFIhopoP9jzo4+0bKwN/ckKnMIHk08MSgV2taq+X/M4XP5ihGkr3O9NEnFDTNL/FZutOz+F2LWP
PvBuW25fuJVJgPyShKUkmJJxn9fIY3M+d8RXdU5L6VSXOmPMu2tr1wMMYKJrpULnmR5QDP6Gxm/A
2rz2R7cLCQWW0T9ratFGen23MapHlWS4Ign5v/q94GdF7XgJpb8QX1IJt07rbNuyPLTMfJfQoGsp
XSgo7HqlwKWD0RR+YuWKb9R2kYno1vmRXjcPFp2YLjlYrBlXkPLJielTPp1n67ch9w/achPaC94N
7eSqAmbHRoBazYAoMZSSHVKc+sgFpXjw3P0J/uuSjwKjAZdTSgXm4UuWr0Nz2L7GYM7vJ83W8mw+
fLsz+RP7wtm8HhPJoTXJYZUGIE4dWDiU3rap636jRg1JSDV6BQykfkFYTusXMIF7+BWTdJabvzxg
xlSjLhfUZIxRPy1K9PzCh9VGGIgKgshQKdyiV3Ed60ck2QIzbBAoSfWJhFVH7Gia4Ulw3TvVZsZD
fJwQ1E7U3Tyaxd/S/N+xCOTYE6YM3AVKN5O1IWJW9xx/Ttmzm6TCs8OtCazpSSXmmEHHwd0k528o
gR2dSmZN6Uq99SUpO47adGiJwYkzZwsC5oPVO0NeRYFpuSia5+jj64/FLWnbwBy9Qcv3jZY7NdgN
HZANqLSUfrTY5CcDRwwRa9bPAxg6S12XJFnmBhSoE/xXWv79ylsAAG04LrAzLufbEzpw28Xx1dtc
WvJXB+xyiuvIZ8MAQscGBE/FXB/TeQfIELwEq+dcsdeV0IEHvJawEdWV5BN8NfwCyYzBukKg8Mzq
pOb26F4GyvKI5Z3mIfCRoaJmeWYX8qfSDp9yXEKlp9HjOmeK+u7lDIWfow9xaR3+Wvj9kw0uG3tS
bkUGZd9/5/1yC+zGXMV2AORslzJkWDe4MjVe/ml9KACqdijo8NFUY/uy7a3DoRoKACYe8xIx14j1
spCDJ9lOq1A9E+CUWCpZ5YWqW4zQuS6Bx+9eJlIUwhhtLDyhYrJzZHVXwAotDpE+LdvYqCBDxCns
6l1/Hjh0Lb85qI3L/4eYxtBMFMUQN6PMDmWutCboMiiq3tbmZid0nUxM1GxtNFFCItv/nupvRda7
+Arjmr1EWKg8q17QsrikB3n4Nxxj7UVX9STgkVUpN0ytNNi+WockiqzUeZh6GNClyvpKSjhKPZxa
r9FB3PhsAlj7hGd1vlfhz0hFx8j3cRpYRPACxY4jSm075zpgYQSc6UcwdsldCm9RTJ110EnEKkp3
goi2ejf5NKrRSr3T16k1dl/V2iajDpVTuAnyMNkeLlssrL+IEC67HpxZunhg76DpLeWywITyWQWx
NmOJpx00fqtgH1bSbQnb31m8Yc+mZXiIy5t/auFf61rCbRGkZb3mBuJUhCt2t9IhxGnj/9krIbXP
9LzzvhQQoYHnhxnEW6lzxlWlxfZSCjOzPWHr4PFCW9iZiA6hHZOtSitKg2jft+U+C8Lr31GKxAAK
ijxMDNA90NcZsOsKhWhCjk9lujbhH6xgTCMeqqVwtgQH8TEtieVWqrOmSIqKzmTKcoI4Nw/2dA/Z
OrjylLkC144z3cgKuO9mHfu27OKysmZiRx0oXcJiGrOLKONPnH8pa6sZmGbbK0rJ+pCJNrPyazbk
vMtr5a4ewVcfcJn5ty1atozJityHElUQfNQYU1KHy+rOq5octSYPdV2cAau6NpYKQng3DPJ1aFtv
x4gblBwAE5Ii2uOiQWpKGkR5qac0/Z8Vny63dMDY4fB7Fr0wazqXZuc/Qn6VAInrxBC6pKwh+kgZ
zrY5lFsDLsb3Zhuz2UbLe3kzribN7HLyQ8DZ+M9+sMVnoE+fYIIu4jn30bgqLJgbA9A/W+zlNRps
Z4Zw5oR+xH2DrWzZsSN7rG60DuC8dZOb98oFe0p7Fiw76ftGDCA8jT7eLsR3K4Cnftx3g5NJQh6O
kWwb3OEo1mL16A/6puFBlKbFFg/F+svZnO5eoKheK8UhjG7yBBb9zlrp4xNsSc5xCLxn7ROuU9dF
yXTD/u0eSZRu2x+AF1Bt4OTPFyFQnee53l677gEAiv3N9+ZYmqRnXFachL5lYSnpU5r9cBUg01t7
QpPmYKLzUzndIcBJ+yjGDH5nSeyY1fQAf+3Wr7mi6IG0h+Za61NmKresA1fZiSRs+MEGXZ6z0YUu
0c+LqdEbaP+GYWjF+o2vCJOamwVGqFTMYASQvpoOu01MQc/xXBdQacGOThOfNnKrKWjXbWSUo8bG
N9f2Dkf2g4i36qd6baPwpO6yWFi19s+dbaIusXXb6XMvLIIu6VKAy7DnD6QefOVm3zOQHg3MSNlX
NhnI3N9oV1fgMuBSxUfgLmFiO+wMCvAX//DxipAabNuGNtBQBZ6egFP2dw6HpC2Lx4D5PdFJzGrc
eavRdb7DGj8bwoUcM8mNeTexgojwgPuvqKVM179C/xOkGlWdq5PKHMlMdua/LMRqsDVo0yVSXjt9
W1vAVK7deoj72owHO4XLqt71hFjQgJvExH9uvy/aRi77EZyM0UXtlVuDbd6zdH4s4y8+Tmk8F7Gh
B+rtSrXT4bkM0c4XvRKMjW7DkNGtJ+ndLik6AjEj865wFncGFhbmKoFFFK8ijG6RGEzJC44HO8Qc
pAf51RijPNkTcuLqWSySJ1siVGZ4yanzhsP2mRMR62hqfndaZOgcBsSDQMoAMgSq4aX802co+ksJ
aPlBRVacORo//reTDy/O7jv0MZwM6d/dxQiE1/iywh/3LOmmblPXmIM8dABeW1ioBKz7iyTDEVmY
otPQNpS01RRDEuDe2HJiyTfkBqxmHiaXyfI+BdHt4y9v7f0V7ZJidWuhPBucWFIGFp1x1SRwf6Q7
VcJialk3TCkhw+l5SeDi19lWISEgu306AfvzOhV2R0nu0Ogx9/8KUvRmGB1s+I5jMggqhwL86q8O
wGf3Oj/ORDyQNwNvgAfVFLEW5rY5PX7MMc+3TTxhTxUzsq2g/+ygYfv+Z/GN7KKsGDlGOuiyBtOQ
t6hECv8JjTEC+Tz4I5/uGxZehLrBZ9dTWvGblIfZX85v1YYVKEeOCmvh4Tmm0gLxyg2toor7rqTy
5TalavZ2Xfu+vnL52+rFLwqIyDo3CBjLcDle5k4m4g5v301MJrY0vTO2d8OdZnu26SKLCgDpI9C5
jiJ7IB2WW4nm5UOFPo2ypMVuXVr6S/HeJ6kDOsDRy4gXqIZY5+7ivtswDfPfHx6s0wdZh5yQfra+
TIENeou+n9DA/X7/lb4K2alfvryLxnaWK/K6IPbIgMPtIrQrDIYlb1b+xXVD5awacFGSmXPYP+3V
7dsreL/LtjeBH1e8HpJakNNin8HFZqDKVBCSbdVM2gQOmQKnEGiYCqRwtrRGfddY+bp90LeFZfwi
VXF6FZK9kJj/XXyI+1Z0cBkFNrpuNqf17EJd8e71Oe1XXAqaUtGRSqy51ctRMP4ZVTJdZFWiCfov
VN0x2sty0ZBoZg0Q7C1rywxjS+YpUyHELGtvTROeHSI3AXQnr1b7McgS3lE1xYoKVMYtoenSoC0m
KU549Zbiuliyk4zIVo2KJgIcNaLqt+Ly9k6hHamWwjTdt0rrB3E2PnAnfIdn2W/l9X23LbUI4BNE
irvfwM8tiGhIRg09vGCrFU8kt1r+wOPhtYcrNlcRavEUaI8APZ8Rj/kHDulJ9EiTdMwDVkdryBtG
++MWsBiH3F85re8McDDaA4IbTnIBA4UBhS/Eye4QYW66uJ4vqzho98bJflPMLlAUnB/ejsa9/zDP
YPYwlin7B0DPX8Dik/RPxPEHN/VbmmdTJ5qe+Eb1x7quhJxowlOF6mIdvfmAuXlqlX9+vsM2hodW
Vt/ek7QWtc8pKg7ll8tE/yKUXJ1r75ZCVnlXvfDnAZL4Co4Q/NzAp0+RXa387R7+D3BBvNdff4Vn
3bifYfCmTQ/IOL0ma1LrcrEI0vetLTSAlBqndExLkxn3YHBfmmxDRXXISVi3nIYMDqKhzdb0Fyrx
iDUMCxLrYOi86PRbUVSMj8IK0ajwu5wAdX0kNL3kPnKcnyhVtrhf5zcdROiGjdunUz70ZeXce4i0
9V9UBJkXpInrpNwqwrgurmMAZ2x7eyrSiPluZi2iUeDuJVJZh4pnVB9mqguewFTpEUospSSuWYUq
itIdKnDyKboH4JwSCLqLavMHT0fPUWY/AqKf++FIQcDN/bSMdDhlYiImPujafvtG+386/Kj5RXD7
kVWXGXNy4UFX/DO5g6sME+P/a5MRssc5x7Jc+/Hj9St7dKfVoiYCytxgs9PgiSyqtGZXnCc5EH5A
HkTmS5yDTK6emuX9UVY7H9Wu03X2g6EIxz/JuVGc7uq45I8RI2Xl33xVri82g5dINL6xL/Wsvwh7
ME+0zlaXPRXIg99SnOM/N682le/mGNMcLzUVdLbXpPq7RBFozrxDJP6NRNJm8BOljb2gJQ+uzVod
LofIQrmkBuHsVZ53kQcKXQ/F2b85yrBGIFaljCaubS7Wn5jhmDFteGuYE1LATvGB9Brp7XzVikmK
VPJAnc6DD/t1MRNwoodR1fiThEIke2nN2rf8RElJ+ZoO9TRCeflSHGSo6ENMXDTm2T+bC4XvZ6mv
Ycw07EUj6xuJS0MzG4abU71DmA5FLwc8mexcSYQaul7lyu5TQ5q/X1guCTOw0+epXDIF40XnguSX
PjRF9CH1yUsKqIlhnY3A67Xj1dgE09akBajkakLhpeGR5LcpU+JgdX0dbvOrfvNma5THWlv3Eo2W
IgxB9B+bxik1DrHSk2wPsrFPGYwKHe1yximPdzPEdYgycGt5TAFQ4JwwxBq3CgTYWzdDlan3+saW
VneXGvFAZDclQ4sn+tjq4WJ6aWiJxFTKH25Ox0AwBE9fprDf2x5/KUK5Txp2DS3UpalT0d1Lyq5d
ySBwPhaZZxuX2qPw2CmA+nmYU9tYP6o45zNuI4jQ58jX8UbWtClWjA36NID49GbJUJsRlCmuxJ4m
lXH054EIx4K/70S3R1cxp8dmE/ECNKtxBUwGaDhgWqc0DAj9ZhafwmHjj6sqCsGYnj/67iASEH8V
yTCHvqnRWn+nGp3Va1DXMUQsfcNWyeMQrWVGXph7u2IMWKgF7DtDEoaGfyqTHFLdHieJ8G45v0EE
Ji/ERgoHOZdS1bIP515zOMX2VAr6Ao04HcmkKOu8Eo6MEjyXvaYIs2+S8POPndGhV+MIlA2UKtWl
G7MfjwlHDiKJPsmQEEv1un+oS//39uUQfK8soLS7CzaioNCQvVQdZZ+bY+W4SRwIkYixPzN4PFUc
pt60ND7E8oiz/ZcwieOCZecx7B8xCMhbTZM/mvSybTcwOCbvv3ozVhRwbsBSaoEj+UG/XkU34olL
c4qWf0IVWLAt5c50Ie3N9p/o4rEWsnepaTgfwQXFqaWUIkzCB82/rWcnOAnsdh6qAJXTacVJnAI+
ZUu6/XssWJFl7thk8Y4ft/IOkrLGyKra96rY5MCVeUpnuRblqyCJrc4hdbM39u3tUF705Burwqfl
IC3psSoIq6dTuMoZwhHjxfdhamK+PF1Ko/g9PsEcsPIolynA2Ae5tYopu4Srt5YMN5MW6QQFNecl
mRf229l/2c7tP80Ik1jouzHwmELhO6Czlu0hch3vFD//++x6vUrfG0NCK2pQaY5iNxxP4YJJuiq4
dkSbUc/fN7gYuNQ3Vfl5X4+/pWT9e15orpDvjHCeJmSUka3lMC0x9am9GKCRJF5zzOwdpDqpWVAA
82RXqjiGv0FTnm6qkiepbcefH10V89HvHKDMaP5ou9cLA2uBtdFMgOOdMG9PlWzVNiS2osVjIQSJ
f1y71qJmh6/OE9BJUhQDuqE4Abn41Y5xvdG5xNguyLK2qGBBsiSQsueXKcwGCdEjRv2ggV5lWiWk
O1l3lt4KLHLQJLeIM+C9RFgixkbsrphnRRJUh3fQM2wEctmrwY1oyiND8riD1/Y70n3F26RpB1lu
ohKY0X2gXOUYP8y2foChfUBCWZVRR37lhjRYKX6PjjmCRbcV7hkxdHyjUC3gl6UyA7TQyVsnqu0H
MDwVKYHX9ujmWBzw/HKDyeObY9nwGitAhZTLMfNHLTvSDXlCUbFG4nD08v0NVCKi2Fr6X4S7NVKO
USocLe8EzkyJAWBT6pV3KE/Mcg4wo2oe2/4Af4sCvZKAiKword7B7xi3gr7xYYOmDBD8vRktZ56/
7uNLbu4ocWMtzgpaf7Oh60sKEON+J0iib9gNRq3zH/luTnK23Nk6cKGw26WoSsQPwSJUgYah82Wz
TA1QXzaGZpit7qWLFimE4YqBlHriFb62I683LuhSI0Q9v8ohjrqevcjBm858jzUW3xm21rmxjsJ+
XhBYVM1PA6wOXWmzwSrZQczPqUOgxjaGfx46raOyGdT097W8ycf2Gwwe212zITdj3mm4jwZZnIv5
x6YTQzrCjHLNsvQ0Qd5ASUGniDac5Ei6WPFJ1wk9J+Ws76R19od3JLI73asQmQw9ELCRBL1cNmSw
93Y5IrNQhClhnVMyU3PmaDxx2gJiDOd2yEdp956jjctlbrd8FoO39+hQkEjXVG1KwrnC7jnLQ6/Y
7Yz9zEUnZZMnpjqS1Gqq+ZcwJoqXGyXx+LBPVuToC0MOx1GSbKivWe7tWfnX1Awo/8gDsd3EW5gz
TbuL7Ue+LBTxR+o5inmmgKHXXpMkE2z8EH2B0awSgpik92nz7RABWRDRRtNeZjeud7VkSW+j8IqZ
oZJXsinOKLem/qmYJa10kOX1mUsjXT4Ttd2xHKIB9VeYDcmisRpOgYo2W80hugIvZY74xmEymuxC
22tgTygjVCJb+9wDkvq8YveaRfCB3lghQQ9GD59ROWbvHsgy6E9q5g1cBfnBnZg2HsLtPrshnaTM
UfpyfzaTAwWD92TxDCOWkpSImra46g57fwvwaf/JUa3tC2OQUmnXmB5WIo+HGOqMrUu1vcP7uW0G
eeQpXs2UQ4mezgbgBGc8jw/+FS6lIpE7l/r6b+ZNPflt/i1wS9eNHlodFVnZFul56irByUdj3q7N
nHICm5w4zCxUC6r3jFO7ioO6Z6ybC+2ipFhw1tBiLW7Ixo+0R5EY0QqKNw+FjDqpTzhlKZ+SkNzc
dGCSkHXHueXJIuKsIZHbw4VPvJ01gWVF3+eKX27klyHUQEXNOc7EgZd2vdHvHQdT4v43glwELqoL
pXoExtxYRrZst6b1iyNrypjMZFzmewRQvvnInclUZ8wNoWhTnxnTxKmhvohdt7hsWx3EtRpGQm9b
kkyRihoKmu9BZzeLypmGhQi0vAdxmoGED59YyCVuAShRQzBUflROKXAKRPExBa8XSu18d5UKtlcZ
D4HaEtSE2mWAcVCAdMPZmZUHiEY9twEwZMwBtE275pjGic5O0FaNNIU72owab5St/XZEjN894n0C
lHTnESAebPC1mMEHz9uM9NPftIbiY+V2HXu8vaGlibx1+61BX3x9upMIpRDjr6TK7DuhG0G35T+e
TdN4iDTkZNuBkMCVtwalb2Z9VIL6AJpwqvkCeTi2sspyWLduqH85uTo0gc1PohBG8/IG/BJx6Shz
ZVKE3zFbS+yqecyta7kLijt/bGV5YRMFWeutn/nyc+qLKltyPQc0O7wS+wWVkRawytgYRfGOTiYn
7PiUi9C2yTFPao/Fmma9I8/c0Hpjg9wyv54FURMx4b1kZ+cBC/kMY+0IqUWG8QKuhBgJ/aO8lLaa
NIIypm4W8ZKW8WkHJqV8HM/vH3NZf7cmq4A8ZS2kyT993IPKvfmN20P1Tu4F48nxrjTixk/6vXWS
wH2mypfUKa2laTMfpVkj0i9UxDIsbkOJuDf3ru6914plZpx6StCzRlvsIix0q27MaSjBKsfKNFog
hNtuBEvq26z9qdaub+oaVrC0R0lpQIKQNja7k+64PDZYIKizhj4vU4GqXEqE0FE4zWMFDseMoudi
JsVuGPx0JVuXAc32867izZm0B+nP8RbOspy4DKFfujUk285qEjCxuxU+NCkpYGkfGmv6h24KAnf/
F6KsiPyOpSXI1/mlU0SdmgsoF4bjo9GLKsTssy71zJpJv/dDqa2+USTfA+I2gKifo7Qh/VzDeaIa
SmKjR5fUM70UNT/LI4r/IrZ5kw/6EDeydKdlv4qu6tuKByrZ5KUlWWZLOH2xJujHjldM93kya0I0
WTGmgQrFD8RAx9FdxOEZNVsCpCRgZGTK8SpUwBMLElBKAEB2RAX0Uq9y3KOzazG0/2MEIZZebZCa
fTIF/OW+K+EIAgD1TbCUBeT4cscHg2VugIYXNo1dOCpVWe8Yyon3jqX1VuVZj/zJlJ5awXI2WRsL
XTwt0YxMpj/7E54M62YbIGMUemh7jHB62GOSxYjlgp0zal0/qRGneTvMWuLOS3arfPUfmgnNtYZp
uD2wt5e5rDWwpiO4RnA1rOGOXgX4dNBZkPta7yhrWw9JY3XAgnJupkFXCY8Xdp+bCucSYHLodXdy
w4Hz3JuNkE5eoqFAzK94Adt/aLrRzOe1MHjyav4+8f3EQAUHfFNuENZ2632bUnhtAYse3JqTYswl
UJnsWB1NYnaSfaoC+MS88eeLY/+qyRuPYDYh5uU8iviALp+lxPzhVt79x9GpZx6EquzdB9lUueIV
aaakdnhlFNHv2KHW+NYi2ru8z85Pgrmbg1NcmwwWARYhP0M8CK/POIKlQEEsgXpvHmvZcd/W2p16
2+NCf8ZFcMX4tkF4X739NfFR9k5S/XShbHQf1MP6yHd88BMlyt9Aw/zGsR2Pon5/FH4YqP3Es1Mm
KtRZYzr5uFkpU1nJ6OmHM1AUaFQ4nTXWT0tn2L/cG60B/g0RRjX1w3WDfZNBTmJ39/ZJbPZzaOBO
YY4f1f3wX0G8VuYKSe9A/c2sFs0Qj9VBYbxCwHcpxnfE6KWdhxtBUoc8t1hEEsOVEbt14W2pMARB
DSDu6Pu6hRAraN467qRbsu2rKXnz+pDRuouv1FTumZ1PJIKGsjmSmahr3utHc7l/HmfP/E1WAECs
AE92kKz4RIqW3x895H6OvR1irOrLfBXJd+e+xQT3v7oijvy6DVyc116NIcGCw6bxrkC8gugWFnu3
x1obtEnSWhTKDMwRgLAg9ZMXm463jMOZP6ZE+kG+nQGPKxiEqTwp1VBEP8TDcBPXnp5d8tvAYt0S
bpn4ugc3XPLoaYJYcgIqF5cIQ3X/FNlx1L6Ycwc78CaB+Y7wMOh8J93Ms19cPDSkRQ0d1enlKeIx
wRfwG0fVAh8pIsp+f/OGUGj5RAHVsEVrBYJA25ckYOvRHhYkurWQZQbaDzTuNjknqPXscXZiaBTa
fqt5/CXoNbGBC+Okk6n8wdBCyUtMOxJrbVfRupHw9OT/8CiIW8lm7XirHCWh7rF2RAZq2qquBVf3
WgzWWccZ61lUTBtmHEUcIBkYx8l5Wql+tPs4kFyMl5hbdC2/CNpOAIeTbW/AYHm1BV2WIljzY9cI
J4Blyhe98koO7vLnUhr7108vaeamO6t4DYKPtt6DtU+7kQLAREABpG3LGWxPSJ0NkImfmUf9ag3e
LeN9Nb7E+RUsqSDt3ndHMaSTwqaCaqFSNZQUpiH4cJIJgpUu5+wW7dByCyEk4BLPzB+rjerGY8DU
j7QsnQwi7OMZCV4/Bed8ki8nh1ZLPUU4oa9HTL5fsqtVd0RZmlmv3ri91YPuk1RAPengNEOgqJEq
xHUC4+gj4t/Uqm8XYL2qgjfHciKlPvg6jpfi4Kh3EqO5hsFTdqlsfNyAb3iitsZkTKuoyxEVT90L
GDKAaIgxteky9j5psA5WMF7tZxUb57QTm97K3V3VjCbnHYe/SZBgdAEglLKHd4cDj6KjFZYh7A7U
FRpDojoqsqf9qotAqFZ0E9RsW2T/gHbZjqtLlURolUBPuvUpiYMy23Uc2o9slgsevhIK78NulRfG
YE3zyJceY6+4eb9JGWHQSiTo0Ht9ExkMt6lxgsH9YledNZahEnrSTK7M0JdkJ4uzGJeHRGzyH0A0
ZYQe+EdIiQwavk1YPbDC87BSBjt9uBbaMsyhky+hSmjeWhYw2t1BVsNfng2ItAQgFKwzGGlcnYLn
W48By9vL3OKR9KZie0Fqs1uYdvu2evhuB59PmJKKo4Zkatrn3j6CqtdlJAHAlCUv31DfTpF6DkGP
udAi1cL5rLbCYYgNUOEYL/8GSVCTZTKQ51hWi4+FM7Aqn/hzHpXFDx4Vo5baRjLaUCBzjktanJ6X
MaWKk31nJOAqg/Z2KWsj8FdlWU3QUe1Gs+1XUveKH13M3o7r2OizN1Am3xArQuo91N4lZcTi8eVy
BFchEZpQ2KpE9I9a5tm0ombyFSqNKhec8WuiadHdlWrx5OMMdWzPrY4sSOshk9VrbQWjlTT+WMJn
XczRluxRjRsgiaiRniE/1Y/W1FgGWlAQ+5RbsqD/r3oOPWgRes0dyQI5+TlMyhYO83unafH4srH/
4Bw7zstL5IH60KXZszp3vIC+PTb5lTZzuRoJOUiJ6iKGnO3CSk/c3dAPqAzyPUnjSuqiQYwTbC4N
221p6PFeY10ZZlpqqu2EEokztyc0O6GNq+bqffAWPsR3SBsSPN8X1VYASePyMy8aeWeATFDox2pV
U6CPN6Gels+mEvUA48pbnwZVI/WcFtcsQhGLkoiL2Bn+pjAf6QdRXOiJJJUsLZ3m7626DaacEeoZ
hWPELWhA82lhLs71xHTLuM5XS5HbaDT4IHTikgXmu9+BZZrmINYsYqp9gl6JGz9udLubD74tCEHh
m6cW8ZoMt9enqQ2r2avyPcrXhFvDPTTE/gf5XmGR0HhO8p8wCwVVVkSSs3HQxbQvBOlBnS8yccZw
RT3t2akfgZm9YaHrZmlwQsAXIk19ZMszes4/sYb7SL4SRk33yp2qWqqcvN0tvO5aEr2xmfgNk/YM
f3p9FDjXUEcTAg3vxN2kgCslNX+ou35LsuzdZcAFfi43Botby/qc5ae4R22jWGvHFjFN8O8mGhD4
S+eDo/zFCrn67sblCtNPPTHfu1D9/iPsYIQ/fB7H2ztXl4R9xVB20AG3/k+MiHkT4twqrDtEVxaW
sdnHiCnfNovdCYgbPLft0xMkZut9VyvGATROuSREkCGp6Oob/OExile6whYt4fkGtlXJVttEXszz
dJHM9JXQGK4COXLG3zFJBgkNPU910RIfI30bG4IgDYPCaIreYW05SxBJVkzdSyN9x9xzNxK7oNlU
B/hzsLVDNOPmGey9gjUmhpA4YmqNU9TZTVty0e3lFf+SiFH9o4Q0pwkrlVgf4CIqAJOP0fosyque
v1lmYt2RaN7x0jjtN+71tbpM48E65N7NlEPTMzzju1iHT9HSjS8fSbry5fuCJjNjjXRfkUdfjH76
GfxoRpR8Smetzwz8PQD5eIdg4PjeGBgPxwoVLvYtuxFvtpnw6G/JX+Tz8Rc1VlKxjurk8gKS7irB
6/MHzThsBV2xRS1ojcyZMteAjm8JxUBZX7nYJSdYWoZK2/xpPZKdKZjujCSPzeZAOpDN4LrudV1y
sjt+nSIosxd5Ggoamjzf1pwQDtEIum0OLLoGD53lns1fQ1A47RuL1UWuqXx5tfd4iDp814yyaI1Q
UerUQJm2D9DIHgphZf4hXwFDzLgy9gk7pikQbisWx3NPVXbXFxH4DHmK/JeKTHn3/fk/yaq5IBfk
sEkM0JsRSn9D4BuPBXuLqh80jZ+bl32aktA7nObdNDVt5hFXitWtrCluZlFfFGl1WLkNIKaUggAv
/trXEzfXx/vBo0c6MyjjV/kvYhmReHBYdrUvYNZ75jMhicrJLXxtQDWge3RJHWScGjaD277aFHkY
qBQxV1C6W3KjabgrEM27Ihj9m+sUGr6P5J5lQiTsMxI5F/B33Sfc4wOKQBBXhcAhCoKpvHgvD1h/
JoqWVIs/XmO1p34mw94zzIbZtNzSSHtvLP8Jw5sT976BRwL6NFImvtxpl1ofVzHoAjsJtylWuG2R
J8xvSXqajXU0P/KpgXn+Jrfvu+Bq1k5axqnRsXZeNzQBQm+EbCDbwUZQ0sAHrTCBLCW9dkmrvjyX
CxPpBEqmEiGDW0QSIiB5zzqliC/rqi04lXiKa671I3tXuVlGoMq7PIlAU5ztrL3iR6m+6rP1sLlM
Y04tRbyQ+kX6GYQKL7jEx10+KEOttPxQPvHCbVdACmLh5rfhdM6f6kkM+0SGEoT7oaqrUb4IeZny
P42B2EtFM/Ko975wpiCB9HaXnQlj4VBzsGKzDJFyQOi2JPiyCxC1WlfCf6ZGB7+N/2ZfNcJX0Kr0
ntaHhjvI6rlBfql9fBPAyzpKc5CM+i48IGtRsvRZGjZqTVWxz+h+pWaIWYdaD2xISbAvN0IDFGqR
TdkFwlj/SDk99lBq8Uh81BKYzKm0wyLs62Tp39TWDyA39zykBbiynxURUr4K/7o7fn+23RzfIjZD
M/vC0LeyiOSeRSf/01M1lFQW0Ch+oHiSqV5kRzJi2JEc2v60VmWwAwT3fZq7rDKcnr8GdKprw7Xr
kLrxWk7VpNfrO9oiDaQIthRgW2GwlWwZzYm1ucgx2LLDhVEBSOfxv/1JIhsNmYYogeyFVNlLPSAH
/+s9isiAY++O/5XP99dLwYLcFvZrtCRR9HcCWPjYMdd04ul61NVwpoVYm006S8wKY+nM7ZJbAY5t
sbzTvxzeR8gJv6AusT1tOnhEj2M6WXesFe87H0DEvYqviWtSCAs9KK9JDCBA+4BsVi8GgIDukCrc
RHEUL4a8mLCA9aCZjxehkKKZUiCRVLoRMhIycSk934U1cYO3kJG3E3TgmgShc0Ea42ab53MNQ0Gy
gKEGRk2HVTEF+JsaEGQIINXQMrUIsXuptA/+6AZAp6uhruu/NrEOHFce1UP14+Qnw2r3U9fzsUEF
qxZLL8AFDWkI7vGqo+znxT0Iq4zW1RKQgjz2cmetRgr6uhDzm3LtE9DnDERrviOosq/HH/rpL2mM
jI9NssRQS509Pr2Cg3ah36oacnXqCSCMoPtySi1pdiof+5U61v8kVmyHQMuzYMX9JlPbbYLChyDD
ziiCMWooqbFDB0LGAt9Oo08SSorJhoB+XKYpDlJMFEiSz6xpv+mTVDWrEjGebW7CzkmdOkgqPNrr
eCBXKsh46b6R7zShvr560JwOZmlq+9QPVB216g32yWmaZO34NnRWQrlCAyCtJy0I2d6HxRmFSc8U
Ouv0bPMNjC9AwImCwf36mi2WssHzla30KC1e2q2fnJsZl7+3kopyOd5Rg8dxrlb+UANcRgubg45r
AUoHP8RG0FXb2nrcWVuwni03i+XlGuhbiXWhNmaT7fOkqm/6rGXB18IDTAWdL217wpy0W9Nmf1uK
xF0MbhJ7EqNyZsueTCo1vPbOZeW9fC7V6Gdnhck40GbFJJ1RPAI6VH6corpir5IiSkcrQpqLmcu/
m0OrrUIO6R//UaxsFn44gNFYtxhW4yrcGBDbDifHx7zpwUFir9tVCUr7qlL9A730h/snnNUTJnam
hRsbUvvtPfaG3KhT0M1nVB8W4JN1q3PLiqwyEqgt+nxpZ3L4wKNBjSygCUE6pCZaM2KcAytzCQ1I
hw1gLjy2ceikkVNd3R9vTbC6yJ6NGI5lk6b9zWxZDPr827fJ9Or6Lui12WI27cY9DzTAAXVQRXwE
h534Djovb8qJ1qOBhL8oY8iE/cDfqi49miovgiUcn4XjGVIPEEKLnb0JoBVprQhd+Tlmo8n7azNf
gECxPLUtizSxTXuIhT7Eycag6Haa+yFyzc/ddmh193H+VivLyI/IXwnPoFujOtda5dk1IRy9lbBy
mZw23JmfaJjoFq4kolJNe/4ZwPyUOozcxOLmxi9pupfNW58bTGUwVLIqUdhXLUvUhVTCvYJ4DEgA
4JMTi95cYLnkzpr6MkOXAvPbjFc7tHoO1o1UCRH0M95ovKdrmM1dIJ/QCHb/f/W1MJkNyYpEe0Ny
vbMDoI1CXm1mDIEBtsmQA+rVMI+5ObOFOuGLiXFLglK9CbU6OT0l6oEoOJAATezMxTH4CqysPsUZ
7I6LJFV7pMnhlF/YGiP/hheHuaXoETUCQ5yejKQvwH3OuoBvQ0VwiaTlQ9AqzSO5GU7wLuZVtaNA
N2eRG/UzmAFcgw5G2tm/ILWA+wKSDo1QkPg4GdSZgWq6z4GBzPqmbDFJswJeGd2yA1ND5q0iPf90
vBVAPCgD3FoYX/6FZvnymSW1TF5iRmaqdISWh7xnOn7aND4q2U410PjgZgbfyB+1MAcbqXq8sIGe
NVxGD89XMC+3qzUiNTPrBaZz3z1bztaSm2K51VGV4dY5awXSCHTj60MFYchcZqaCXUp8wvxZf43v
EaS/glwyTBNc8PBLX5UwRl6mxYDW/9QBkmxT5AHSavfm5KnnwtoB7Sx5SHFFIjvXAp5JDt5yqP/m
3nQPW3v7BFV2E3HnFPzwRUpqqTkb0GN7D3dSgSwzjfe3xcX0JZXlf7oXLOT2fCaFPrV29NxL5Bdk
Ftx9km+r4wWGAkv6FtpjKhpgEctDi0fIzQ/CiMWE+40RIyMX2i3+VR2dcg20TV+fytbG8sZy0c30
gX6PvCbDKZlMCyMo4Kom+HDdY/ElPACxPS4T5LxfxGWNXh+JbWjsmWJyR0uLNg+PUeVmsZscY/XD
buZ8C3z4CJF7M4hvEW/3eUem3s0io/Oe+FMdkuBJtSOzxB0ZXAhJKMh3coZaqjm+LTw6HM/djoof
0kp2b7C7i2y018GrnJqVBGh9NkGWxo63cku8Nj8apvsx6VBP2PRR0ApjU+4VJ2Eh4ASSm5wJVlOZ
IyOMqyHA4wiWr6Ce8Ca3/1X2vMvg3qZ1qP24q3hVWNIMXWxqWPvq3bSgiRmmOXwnU41V+6fvYKT7
EHaLDD8pKyKZ4+rN8L3jtI0kR9i/ffvC0JunsxAhRHceGxTcHum3Ru8csFqkE7qRgLs/FV4bMsy1
hME8CUtP6BGxh6HvvlpO4aROdTO7tAVVhA93okrxNRrYtoKbIN2IMm/wwNBnWfgqwpmYFD/2c+IF
XQvt1VjGgP/EdSWsQSjl0o7N4iiP/7UR2qYJ3UDQaZ+YHYt0NJRVb5U3ADUFxKVkQERqIj6Wll17
IrtpACiCJRcyXM7n1v6fqXb/poch+nKd7qNna3iBcAAdpH3RKuEmBVyKuYUYyMkdL6E0FOwBeSEK
aMKKqWWEA63thcXHT55OXpiw37ElGX1DY9hT3a1SqcOs9DKFO4EDkwCIgAhwXDRzwIgbMc9ICNad
xlwk7DLpzEsxVd0bhEY2vurY8omthSwEh0VdXP7pUGyGtprcLgMC6SbwNZF3l28zMSAHyjiD+9AG
HP6P/gwsEJMBQ3YiwCF88fGS1Fll32ROGFreOwUJ1cpS0k9GIAe2+Os8IeOjQpnhQ8rVXnLTnf0Y
O0RLxUDwm5JBHS6OxsvHqrWPiuwDL6l6az/3UWJIm4bza/PwdkSzh2BJNjayTFtnDP/S6pgkPSbN
bqlu0+B4Yywn4J34kjMy62zk1/A+4Jh1fLM7oQWLNmonMP4G4zl1DGtXRmSI7TrJF7k1bNu4YUcj
HuKmHI9co231cJHWYB8dB43fNU9q2luRAR0bGa96GqzAFprqJZtmVR568Q0o8BHSxJT4eGY8V8fI
CUuIy1NszwSjfKGpli58eybtT1tuxu41UckSQgz00cKS1pDxuYu8fvj6oqBIUvzm5ufJs1kUNuUl
iubpbMm5XyaSGlnEz9XNFYnPJBKbBWKIrzIObrD2LVtkTI+By27VxNFsEM3j7dabiOUdM4C8+oWq
KmRaWsXElH5uZbaoin4mxQksADuHqmDMcl2mqv5GABZsoIh7i/zTbywATNDZVyL0mkCCqLyof1xh
iyRSjGGmBjI+MHI6NkEhKuKL+ruOSm0VGR7QF0jPU7w1H1BO8+6mgPqjKr20HRwY3v9ADa0SAGhg
uTKsdqa4HbflKFRHOf4MsiQsSMZEnJCCDCm3bA6NmCgiuiC/rIqpeL2qWWVIVXyDCqp+9HFvQK7o
JOseXnpUBs+XVoPVF0YkKeGSTKUy/JlMZKcMwClsYUSmrreGvOw8RTGkv6J+aDFXRbz+H9VhBRqm
mYIq3gFaZIaMzxEDqYRoOmgonqrTSFHDNhms3DhA/3+HLbQ83aivZg7NuIk8ll5LnaUi6TgnIx8R
SFP8ji/Fer5KMgsPbWM5bmSmTqt9MDzb4xQZTWvDBcUUKSVgAk6ChCkRYdyFIA/mzWqaqtdr6t/g
x51+WEFHo3z8iCdo2rLrHnKjIESHS/+2c4+2XcLaizS/FwzYHrJJXFMNLVsUth75eO1fjyeX5HFE
KzYeY0J8xtvS4m3j+YtkIA+YZ6oUVr1smJCSODVlgGruIUg+vJWEFQ+WCROWx8S1GfUj+Bg8bFxr
vChB7gyPg3kLO4x/+f0Pzb7CEhLSoa4l2B6aGneQYWxaMMDrg66mTieqFYSmdgit15ZBJgiYGubW
615G4g/SBsKjRH8YfhiDZmgFrbZBOyCSKvhOP5KRCwkCR1rTqyjI22783SKGWH4nwEnB94jTSHSB
xCIjLmorH556JTXQrizOeMBjFOOwqofL+WrTzySNFjW0xn6z/+a56fvHNV13VEUm8af/j7fWFCsX
dqNHysqmuBKS5qfzmiwjHIcpbvTkVX2tmKduDFF4OHSNdshz/sUc7gHlzcjw9Mh5o/O0EuPb+Ip2
ull8Cr4MN92tpVnXkwfls11LizdVQstVOXo6Am0BNs9JjO57joH4D7q8/RWpvdjtMrubHeJtzrVm
KVRUWRSYGHaweUQPhgBqWEAz9MZ9F+hrd3Jl4gnH0iobwimO5vNGwamh5I4JGuR+xWXzsXtJx/r4
kdauAjwktfjw+oIYT+ihdHlhV414ghSa0n93J0vf/7jExoFujXG3V0aNbCeulTBJ5qp83Phs4m48
KsULb6VrXKFedArhZpTKpTZqrFzyQhMs3vAWdrJdCACEF2hS39wG4O++Osbn3k0Z+/kJzn5boGkQ
lZRtydwLYIZcH0acehha7dtVDbSPsgzJqjFEkB4p1ja6cP/DdXAsqNAM68tL7ITObfAHzj9e5Ma6
hzvc3kV8NbvR28GN85FHCNzlsMZdarbyRXzQ64SoVmWblxPpC321HeIABoWSAUe0fSG0UL2kbNaz
jNY7qvEPB2YoYYds7VPeYydPLsz/e68fwPB4aiepUi3YrFRTETjy+bXqtsmuaOJJDgQKcQ5niDTd
Zn5x5BH4WPUCwVTLSbpofgmXY7Am7whjFF6yM/p6s5RFxp6RWvWjboBofgortaCxs2/Qy1PUtV0u
WPaxeGf8RP5tE7IQmxJI02yKkGkgJXR4FO3KFn1S37HA/uCTlN8UM5KGG9yYow9yeIVicPEsVe4D
bzzg84hm8eAMgqpYHax/DxQclirjAfHcMnhfvZGDuk+4yenxcjO30ZYjA48Y2tKTLEqHw0OQn4As
j7iToIMovheUZdGJ3SKsAAm/WJLTUZ3UYfMqjY7czSs8Ta2qS8gOqSqpU4Xg7KYjQk2eudsDlKVf
9rnqFvpsncXjB+1J9EGTZMJXdOFHngHpK6B5Av0lKGF7UR/8+1ePfqXEVF1cJGeMF4H0OAsmMj4U
ynu2xyWbaMFWhUVVkfmEQ018LJCWmga7h6OAQczRr3ztKQLswXflzjz4RUpeew/e3aWil7C7YQ+y
Rl87NIPLujxBnfYY3TXkcyoigvgifwX94956Lfg/5UVNSWGDSNbA0y6k8OwYJ5ufuV/dKiwdTtgb
/n6EHiYf4DuKOUvSBJZxT5NBh17ZdioIV3eTcQjaJRHDeKoeQlNsjGPuLwnc1PSo1P6bqcnevwmf
d5CMZP+rppU5clK1b/cTzt3UbFpQIkw6kAf6nlo8w8kKuiI9kofALWILu6fHifcONvSXLAwyPg10
fjCO/Eifc868OcowzdDez5gkwZtyFxP8Lo6IQaeVlORidPziBw2Q7XXreiaXUAEW5D9f4EadcY0a
Qt/oF4z0LiKyIuMQOoyML0PAuefwbCSokW9bSo0ENEXIk/1+VkfHaPEn6xoOhaLA2bixBI4NcVFt
by5hlwfglImISa0RTrPEvD/vrCiz6OO4neHGFm/xRtXa6gsA8oBnoUjDs/7BIdJvJ05JdlbAn8Uc
YxF6UxboUJxqBonHUycNVzLq3q32u+q7wefn1qTV3Ox0t/TPZlKwRJpOoAfFzPhnk7qGeBGU+RhY
rDHx3FeBaKqjhjzXIvK/yF33zC7s0Nfq6dxbBE3qRlR8j6kbCXxyrzx9trpE9WNp7j4Cb2HhFyNA
aavaDpgRb0DElhzbYHyf3YEvHoSVc3QRuaLMJSNYdUVsHGF66sueH467fvixolmqN5gz8aPy93Ic
EqzJpO2E/WMvY9mJzrCVWWKEFKkXz6mrnMQXtLW4TRUoIrfsEvlWleh34+bpBckxbukuBX44iNDD
2eG5YaN/Nc6Sx4y0/yqZfTnuXlCsiJeOZEZs/AcuEoqfxvcwo7pD0Qp0gkK1Y0TXPcYQspkVsFM7
iogPIgK3FXVAZB3yWdST6+8liIgpq3m/phea2LTv/m1baOVuG5gyM7jYz/PFRQLX4epSQgSKN7tJ
k2IlK1Fvn0a/l5fLrgnle4fI058B2EkwXTWKuiRoDFSZ6no3bxe1kg05gjk/cxL4Bw6hinPwOpmm
Eo1muzAj3uZ8qPVkXudiHxGJQ5uvamfOrvd2Ry8ONYLajw51eqQR7017QITbIyMEdeANk0uarNVW
mA8fB6G0vFT++ecRQXstHos3+4YzpqkQbMBQAoUC/oPwfcnAz0JGWqdBTNflKRSxWELNYR3dJSx/
KDBDT3d7lsZbyivT1x4zj7kOJ1wA86GLBV/gr/fVkAOMB0tUEbBYLbEivNQTTIVsOtu7hvR9GcEE
F47k7Y3HzH5KfRjJet/ELrm6n1vOqwD57nTpPttZeqkR4mKLfuTo2B0a2pR1aIVjI7EJn//lqe+r
NTGKASJ/6QtPxlayfUOp2nCx48qRfFPWujUjTRjVSaucrbJDtWHHjn7DuJlyolSaLmcEUh31t4DZ
xMb7/mHhcfxW7zm2HSQi91R4TDn/NioTABPyk2lcmOaEM2D3IDcuwgX7StAzclzlRI//hMrA2hIb
fg+6NcmzGKZvMtJKdIwb077SH+HNH3jV/gjBrtQi6CCiHw2USbSZolfVoa5RBmMw0czEwXImsPoN
jOHiIYX+FHGvywHdEps9e7RzUjrhlHFhIsDIzrO5+Pr+6lTPNkOzakFHZLx/B6KuxVROru36gYVD
aYdARnVJa82zjIGeGub4C8lsZA/26LzwHDF/Td8wUZSRqiUpp10LNE5ZqL4K19ER7CdbVUwQTf/p
EGa6Y7dL5zb7S4/GK8VchtKZjOtL7KyLDhRCboAoojZ4eecCQNvafuyanjeuTo8lGEWR99H9rbj7
k710wxZCfHBHombcsN6tVZqq7Cl1hapbMlYaNWTAIgCMMAhsOIlDWLmGr8N3AJjrR4824k/8KmlN
td/JXhJIov+kj6EPhJRnlGyfqf84NvcVxZ/pI08VDgp8fQwdA+5xYd4wZFK2/2enW2DDuGmiS/3H
o0eqF/vPH97hEmWvwcGOCqFDXxmBzOz7Y/CV2pVNqMH9Rq6SY87Zah+UUFh/t3mzoZi5OzIb8gxg
7UInxmQn+KTqTrfPmpqUrC665eRMRCU7QoIuSGXMyIJ0is1YifZAFgriTPJjin4aVEhxvYQrD1aI
SGRnzKtPENwLU6DyeHcLUnVLCk+RIsnxPcC+ohqFH8MMILcK3AQSe0sxAV5Lj2LLMpp7WjKZsznH
wkyCyk3wvH7pZn+OtfRKQpbfxFouR36p8KO1FifTLxH/2cqybPtnrNjOCsrvZJueESvzZj88tCxM
oyyMC25Rxu7YOeILtwagETVsBiT/A7Mh+Ud/ctMnEnvr+YbUN5iHslyBGxwnh3WI4PIr32R7QUEX
oRsayWOjbuzJkbggvlERZSYAw/3cULnfRBcVe0T+IvGSCO04vi8ypZ5wJ9t4CtojWkRHFfKRK/Rm
aY2PNMWKDdqB1MifqUyuZGc0YQ3gy4jz0jM/sPwlfUgXIcxZS+vOAddmqCXbZkkMO5VIc0I0AXRa
4PQv3Udf3F2v6dbmb4xvUeWBxriHiet1VDS/zp/7oRu0f9T8pJ18PkPj76R+F8l5uLYp2AxHaC5U
a2ELagnac7u6RfAEhZj/C5b+G2xVOifqOaixJ5/fl4GnAP+59lnS9nZanzMo9z32Y9TM2vMhrqXU
Z9w77/KSihPXHzaP2Ge4v4mCa0+WY/wS2sn38/YfAx3U2pl5BrHfMtHepklxkk7Hyg162zPlE6s8
WwXerCcc4YzpNonhtaXsBs5dP5NgA9uYXlB9g5vl6af7xEj3sX/4k8rNw1pUb6w9eoE1493geL40
UO4MuAN5aDKO4qPg4ZVNNaV2L/6V4RVQf/etImJDwBG+XoFS0kOjdhXrYQ8HQyVeZExiwQmCw3tf
lR70k3qtNRQvux+ptJplHmt1CQtqbCjngvkbV15xb2AZtA2YH2Fb/FljiH/ydYZPQg8Fg25BAn0q
m9Lzd5vOH/0kRJn4v+aIb6QrMJL9jVcgtfWri/lOFPvxFa63yzS0cgG1iaZOFS+bQ4ABvb2kXPIt
MpUpFhssQM92tSrCX6ienD0tLBLKWUkytGReMTN9YeZnsmE1kDm2PNwLvcTs3nxshJmFFXgxpyFS
3Lzt3cxFqeijNgU9tEYON90aCVbzjyF7LcE73wEZWoFfNwV7MGoQXZo2FxSCvEh8Z3+eN+ktx17l
cNope6k2MforvkQKsRkVhdQ1w1GUcWCithIUcc0gVuNktyP8tuUwhkkawcL/G9GFkc4r//v6NU03
bLF2kG+RVGBrkiCLPF2XTL7a0HKfY1d+oXgJtVLlFk3cEYffH44NPLfLEZgaXBMd2EGjFWGXhDgK
6Jnm40BeEomTcgO3gW4SlSlI7qvFBVRR2js3xsxmprfV8kNdwztO95exvWUScB766Y+uoMIURvlE
qg8Uy0EdC15efNPnPGNKjbKscwZ0v7Sato5dPIYozQOCVxxpZ9JcIsUFW0ITMaL8WBAj9DL6D0JZ
zlevEw5KUNk5wL1B/nUO65pgchCpbgawWf0K+2l5VbLSgxbs4PODyd7C9rK5yqKgkCnigI0js9+X
QOYAYEG2fbDj1tdFdkEJIxkN97FtC8Bt5PWhdIELUnfflwaCU8+90MBuiRTXESvloDKLZ9yO7DaV
RNXfCX0om0IU447HajCDcco8ck/E3eNVBoHzMWm4eLynuDXNZrubQTKGMIrSw+U3ZP9nIRoRVw4J
oVcP7T3XbqLzXbXnlciIyqn4eJnJ3tiOzRktTMUsw1HEYbkekY0YCEnJ4l+pb4Sv94ahLzyr69Iv
P8n70LImLjBUj+EvC8XPllmr0f8ViWmANErBSfAMkH3qb6nCTuEOcJBM2PHbhugW/tVcPaMARfwH
wJvL8Ha03nvGBubMxRRdQ6bBZUfS9PRKBEeN2MH5NfFHE6+vLtyLrHp7T059z65ajPKDX+h4gerw
93jMBLEBZ7nWaGfEI+QofjIWxMIDr5DlMgcX2BlWqzrTCIRF8fYYGBXbQY0FGqtoa7qjCi+AdRJv
FJPT0jRs/6QZd+m0Bt+uEPIVXz0+HlKKMa10siynuE5hv8OAp+jPinkYmH3h0DgrJVgfUUYGWYeJ
FNfP91XcDDU/iPLN8uMaHr6GcR5D87EddKEHjDWQSJmpI/neoY3f1ANYE/Psnd8wWyjZz6tTkkNb
bpw9ESuLcQHXZti1a1OmUn8rJt+UVNWgOchWGC2Eqc1rNSjp8EGQrHQxeUB7wLXd1l0NQMsibKWx
0p8x0mWAz3OLQfEbMVq8fxttIb2kulNMXhI9z/xa5kSah1/IIUvfrcil6ru3NCMvh4aKSdUTa7wl
SbwyaEkcjbVIxszrDFaQhSzDj5OeLtIL512KZ6n5K1eSK/d51BJxYBuQ7rlMNHF2GSza/g4sUNFa
yUGtfANDiFc8a/EnQEc0FwlU6JAMLQPTNZsqTkCI8kbn2dPehVYE1u5AEdjhjyktq57UvvJHr9eQ
wHrbIinvzelpJxHKGb+v6LELsXbF98TBT4USPU7oeZHMlPYFiJ5BTiS94u0vjFWaI5K0zOMmo8av
7U+OL44yhpbB422sGjS42ufOb81vgrxtnX6pXrMRInGqVagtFwpVA3pu8/y+cqggSa+xjrhRNUaA
4LGtKwfDRUjOpmWWN3BX7qAEO/V9xCw7FF3OoIZUbLN4M918ZPrNgmXf9XjHhEbG0ZzPgm9Nh418
bgFbZMkGyUFxFoQ9dtCuW5xdq50LsD0rIcNiExnoA/wRsKdPWYcLTYTvxVnHK+uLUIdNeYyUJHMq
ZGgwdMJFJlamYvPeFrZassDEXnoEEknp/B8IzI3iFMXKvV3MpnS6DMIYnL4+KdYFS5csC3Bw6Ita
aBGwS4Fm7AHvrt7oJZWYyUVHlluJVzx5tgwncNneJe1rznHxcFUWOaWUjgkEmYo3DQcaejjic3/k
L7skwURO0QmAnYf6/uvrLf0w2fd+dAXnIRvftNZItb+5rDUBHZbe8cDpE/lZR4q26NOPXfnp9q4j
0CnhvIC4otFMvbAm5onGqlJOmqyH0ScVZo2No+6l7ok4QndTWq9HKyciP6zwy1Dxa9qW+nmitW91
JdegG5FUEDs0WA5dgZryUpJa0CJpwY/mk/T54og3jBo1J6ieaU8Bx2Hw/RQHC3kb/wjm9dHLcI2K
GxsLwfhCl66AabxainQtJgqD9EhcIKoCaFAsr/ZReeDP4MgcYm30M2vkvorAAmwL50D/WdUWeGIV
GogbugYaDZnLdvZG/bGHvqNy/xAZFOxk3Hi06OIEWFzu3cxlXwxu5eoyN5syD4XP3TOmm6uO1M88
rU/R4oDANmSP9B2RXYZ/4YKgrgrwkBgC7LdkpMdzrHmhGkqZ/zA1vTECKIJ93SZC1+Uwsx72hTC5
OmT1TtbrbsGcDxP9hcLPNq7vcbs1c0qsPuZYWCHFjzzA2B0SeGit+tZDUZuEmBTCA7UIeXMPyT8e
7brYEF9tkG0+VZ/JiQrRgZEIhgUzkCNKyAb3OtGv145Qd783t8LHPt3HmZZ02hpAjWV6zx2pspV5
UsEGQkTzr10dSe1pLvBWm53xYz5LKdx2aeUwDz36jtOWRqxwyupWdWQAOF4S7Of8dcUW+k3+ne9k
0O8h/AAWHVg/XW60FulDbMviYNJeG1JEaCHY2qVO3kXqJGwA5//LNKDEU6lXB8BA6e7uPfRuLP4I
t94idYhLn68Qi5sKXLhsH8HAk7nRlX/yGgohXXRxLunx57XJaQeEFRotCFPic/NGib86q0XS5UbZ
J/ViKDsZCvKSq7nx1XTnh+ztF4JXywATXcdfrRB1okbKYcM2ntlDbbVvwT46PJUCRsrMQAmM/NYO
W26aLcHHfuPGa16fUgGYH0yXWJSoPby3IPkosw6mcQ8o1awAm7hiIloyb53OcYezd9aWIw57Qd+l
7buDydYhwUCsaXQbLsUGH5+8Sd24PT9t459dfqcKbv5tSQbGI5Cg44LeIxcUFJU0QF5X+lO07G96
yi/X8Dhop4gm+lyoaFhqczI0IEoC4z6CtG9sCM4wVcORcmwKNssB8GxNQlXtwCiHUx5/VV404A7y
WPwFFrQJVXbbznD1Bv2aLU8SX8akYFNiuyd6fPqJBzr38vSlCEhkf9qXUP3gPp7agN6/n8SQ6/Vg
pS59Rgts0w4pA8OAYVEyTW08ne58nXwrWEW/db1JNCrZF3jfpCUb8aWH7NBRcNUXRkvL1YqKCYgr
ZF3ix0IRWq30SFvU72vYXapdrUK8UFXy5q4unVURwDqP9/a1jeyIT1jelQrURMyX6mTnPRqR9DCP
bc7HwJilJFzEVbiq4VLCMj47dm3Tl1bc4hJoA/pjAsSpKf/Tczbdroqm8W3E9GcwjfVURO0Sqziy
23MDAEOfOaT1N6cju2+Xx9xmKyTqGwTNO90E/GUViKCbYVAr9jdi33WYmGrjeci9tmXmXtSPUEyF
WOtRVySoVzGEAS95E9wSXY/iH8Ihvxdpdw8T0QmZFZ5ZPkLDawdTMGNCWwa7/jJ24I4GyZxBf7Wy
erTzpT5HHslIt0V8+mdU4xIYQE9R876iKtfrJ2uAhGESEjgRDcPbQ8hWmNZw34u6j0r9o9sP7dle
gyKm1VmVBi21oHP5D1JfilWQiiFTBUhX7RtM6b6krpuhINcDsEn36iQgz2FUM99Smmnvk6UlKz2n
b/SaHrxLJi0Sj9bfOFep6cPSnmYyCFR36OrGlfgX+CsMH2+8BxpVpZq9vpsi8f7Siw4zDVRUkUqt
KSLZWVCpWwZgIPVBujFYlaivARkRCPYBnJnNaNQ4fYNA7a+DVXFoiu7ubEj6TvkiJWXgbepwWHVG
sm7Gy39nuxYR4+8HbEliqEkmvll0KfoD8z79Ba/O5gsT6YUzniBk/hW45fW34NwG2nmyOky4KWw3
7sMzrt5u+pKG0ro/VITqfWLXh1KmCLP0qCEY6//1gqERp32vk56HzcIa7r/ck1NY5jvRDwU3yrs6
ANl5Em4IP2p4WE4whKaYSWNsLaWVqDtun0M2WtyPjWEApHX54F739JzSizDyxNlX+kZBhWgGE0eb
I98KmPNcloNPBR7k9wjDQmQN/N8IsinYSzcYdldjuLvKbd2Na/olkUgJ6ss+t6i5sULBuNugeVjz
OA2Hpv2x8UJ6H29uuyEPA2Q4jCnA+rYgpOQQEtnu69F5umNVcepOGXLDkmebMZF1hWnwvyy4quLW
6/DlrmaIaqJixvabqmPO9za0bTw4GehnVoVgLPE4SMtX8lPVGKj8XeraRwLGHJ1teDdm69CuEAHO
OkAUt1lLJOX+psD240+oZbimuL71i+/2uA1fGc1oVOhpCrnj6nlaNgYhGOEDg5weYAEQNQ3mXwOM
qgYIPNgt+3WqXaGOOY00BYHeyUTHkde0KkCwrG7d/424auBeaZlgkLwNdEG0gDDbb+IZ7tqjKCEr
RCBK6R7/UjU1xRJRU7hlG+uOpQVjKftxPwnGrCG95T92uk3clLkoZpLFvdCOh1cFSiOWcX0F3fAD
BFHvejwPpEGOAp7cq/+KBBpfGs09KBNF4xNTW8dAeLNnRJQt9Nrl2qZea/DMmjBRVopOUwyyHR0s
2nrIONthbjWTqy4YIdxtAlt+rylZb/JFJd0roUoHnUmYtq9ycNvuhBuj8ZP5tnis7HjMCuua+xR7
rCb/U2E9GOU0poM/O+fHlrsSHMpohA68sL/QCZTUglkeLmcduODUsS83z+UizuSnYkem33f+yB4r
q0+OXXnoZL+qZHEvDfOzdkiRz7puU4Vvk/Pd4ALvOnHQRmE8v69sOnVdTjQRJTj7vN/v/B0Z0mMO
Z9Z4he2l6aS9+KVPBj0J/XcoMyes1wFHKRSmHGylSiwtfBLnTjgdmwVP4vbIvkQpeggThmdxLzpJ
c7NTItPs6DVvdVrI/xNp8Gkm/WCO5hUquFNqONHgZmwVDBMHk8s9vL2pDeJyReT81s40tYC7GYhl
2gtvWPMC0vUztBWvkmzBjjmXAxRkqf54C0iuEFfpOIzroqezCyb0LMWlnkTzgCCC65HcVNw70fPX
xK8IXLNnK3HxvtPF9+0YnwJAu529uNINCdpq6dszmy+2vzLpRIv20k6ECtlBBxoP2ieNrKug6xNi
sZbjCwAosGj9DeVJui5QVuW23FqaB3dDJC0aFkxsOmaqZuXxf6em4nBxofjhsY9qoOA8MyrepppB
WzlGdjTII+ebjyXCPWYOh2vt4OqNq0BLA646oJ/E3c5ac0CI2wC024gltGPq9FEbzVKwUi58nMYY
NL/KZk6Z7jaVAFsEVp3R435HLCskYm40qqa+gkwFUz5kVkIG47qCuhFRKkOuVlXfT3pnWpv+IT9k
Kr21YDVLxc3oUR1ov10iyLtsaR1SlRjAisT2g08kpdds5PRvRVwZVOZPglo/VnWxlt/PBwwJyQ9T
P/josR3J2Kh55UM0E7uROnMfjgVGkdgEoC1zf9HscJZ+sPsysmjV+6AKNgj/3DFqf6a0XnA9fHXN
3YHCGJDwtbO6Z5fnInHjnpkNrz/49yElFy16bB5iBZyOEp/wgXC7wBTd2L18ZqWi0+sUTmpUGNog
eghmP45IOgsuncoyx8vYPfjuLC9MHiGu9IUvI2uQ2QCKuLguOIa3OTW66W9v190CRgZEdCjctOz6
TK2yf/rIOkTLO7aQFLkeUJaIwy7opYnI6HhXT7cNJfxoYQaDBFsC0DQaZhFJ/A637Ohqzl45ScEd
iPJ5oVceY/QzYoxMtuWM6MDzz/7uI6i0LDSyl/s0YZPE81EDr2Zs1peBa+NLZq7weN3SHaw76sXX
9TgkmjhN19bfDGbXM3PR0tkND5ns9t7oyuN9AOUfhJ36oqwtVcHXTcxNTSIld4ZGsx4j/Hm8/sVp
n315AZzGFdPlXxdrcTG7aCG+frGqcEgHy6CfkaomRC0LvikzfkoG6rmXLezB4LA91DL4UPYE8dhQ
1y1RxdKRAx5CiNb88oajvJuExmOCEZnnWcLV000eke1sMbJ7tKuBJ0/Fs5cfkt70hcJcx5sQ0LFW
aYTjl6BOzzfGcdrgwJqOY3+afE0G9t8hYN3TgS4sFEAVTXtG++m4NPkGIG4dtYZESrtqBVJc2oRG
5BJvhD0id7pq+slKIgRs1gigLHi6hGKVeO03VJqcHl0+7NWRNM9L5yulpPGbOV/n6Sq6pCWKFpzY
2Y3ocS54NYwez45ogFypW5fe/ns5hz96XSmP+1nKGRRTptlez89kDi9NZYY4rrj4UmMrn9OV/7Ta
oGRj0L5gsaH4EyzGfaWWoTPE03A+FfZH0DcXDRdkpE3H2SR7kCK9HKQBHxmwsSliFJFKFT8kbP4l
W4/VfYJvmxC8NcMXFsY22mcUhVELAqPBiG8E5AyMUFM6OQ8Zvie5+LmtTZ24fyh88vX4Lf3z4Y80
M7Rb7ajFoHyfOjimoajWO53YoZT5ymnQawV3wQTJhgW+oT1jGHIfVSBbFbjkzvPmhUfhS7ndf/5Q
srs8S1wEJ0OcFAbhhNgPaXnhnZG8QSH+3zUe9l05SS2AvNzOth2M7CzXsWUD9szd2dT4ndVr1qF8
x0n51q+0GBNqMz03peAJUFXcd2MbBSadoLdlwHQA7wpNQ2fEcnHTkBKkbWYQPXO7/RkVDhlyMYNv
aFFE8MAMV4cAOwJw7pMptM6mJq+TzL1tYXWntJJWR6w2usLqS8xv2wY0XcEvWEBQZ2qhlOgje6G+
JJQ68H1Yv7tbC2Cil3zehLCGlmlg9kXZjobtBBxa6KUMZugWkv4OgZWxk288QCpjgC6eE9yrQb3J
fWKJUkrzpky7A3aFs3B77Cjwg6vIZDLrS0JRZaUtifilC1LhvcXsEt7JSkSv8QKo7BzozXmYNUBm
HZk9ju35E58zM2FtkJYJRY/2Jbl4DF47utY2upofj4S0roPdC2bQvbXLePQF5lZt+8hyCkjGZUEa
EhsnryfWzybxe7yBTZx/47EFThWo8gXD4N6ceVQm+bIB2TA9X6MkM9Fa9nHieWNkFaJVczZilF/2
xjewiig/8tqAB8Y+WetHap5q3yOgzMUwxZPNAqMurO5DcyOmRfaDTEZ+7TS/+TlR+vwxxqWHPsk9
ruA3pBgSqhybcQ+wlg+fUXMzvBWUhk6qZSl5A13Yvl/1WNsdWpd4bKRRjm7O5N8n+4eXOwBlm4at
9Za2Nbj5Uv+pd6dwwJ/gNAmNop46wKltV4fGL95o+WHIlV8qmlCqPpxRvrGcVyblF+EvxEFSWD+L
TW7TX/Zi/XQDkM540lAb1gD9yAGfqceVA+5rRZi4mOK8xjLq7OSkL2nc6NX05T08xapAUlUeYDml
mDzxQvnmyxdSmr0eUkevJHI4Zr4keqQPJSv8MJs4F90FBSVfztcS1/M2ivn54eQcYEIoSIG5XIXc
5/5hZMfpt0ZsD7Fk58HKOBnridZXcRD8k9xEcavYAejEyQvUWGm+RpsbCMCdIy01C8j00ySdvkB9
jNm8d/cvvXqvGxagZOxOkhM2gH8aG5317qoBFCKcotORrNpFcY2YGzMcJojEKeOHhl/hfKyH9OeQ
BiC/w08FXxERiovaNtWtJ9xtorOERLNExBk9HDf1YdztVW/Q2KvUji1A4Usk3f0HrzQNwrinUJqJ
bYLIA29eLp/q9rZ+Uuv3ocfi03ExSoC9IEh7DFvjcr6Wja1xFauUTOV2Jevel1y8YoFp9Iu3b43+
8SjMtGiv/3AtlwK5uHAWA0ZkQ5fGB/6H8MwpGs4NaIKqVaC2h3YEhSvP5HV8rLyFIkt+uWunPced
t/n5/4POiAbIL6vVWu1mwkyG+ZJY4kQGoIJqCxb4DBBnRJVSBb5N974UC381B/VXPGJL7IFFTKWS
T5pz1ZqTsx0jPqBDrJNdDoFgLS4WI8EMpnrGTUT3QkUgfpJmkKvsZU1/L2j4/TihbATZObBp7yQ2
9m+jtlbu/IdCIFetxKE3CFoCtmjK1BX3eURNLn/xvF/ExcB3tSdemZVQuQaC1OsxgCbrP86k2FBN
LY7qXrS4C73BYiZlviDaYNBmXlbgAiYIm2VrvF19NeO83S8hYrTQlLS01MMTETYcL0b4jgjKWzuU
Hw2YkfWB6avUMzxFjc1LJKgkMH5gtE9tUDrR+o1fdWT+DqNAGfJa/kh5zK7WDcj1w5NUXf3y1oSc
SzVnNUvW7aGBZokGMC0SMotgotfEVcqoSCd7++MEjKZw0a8STxGMPHOT9/6VYPF1+WR0NcSHGJ7R
Hcf32eWIYRZtiN+vPezObR5PYM0urhm3BFemitFOAW3hE7WpHEuRn4DWiB3SZIGbODkMF9hxrTwW
3h33PTCPUDjR9ja6wdXwvzrvVKfsms0zCbBkK00pT2yRklM5J9Y1lCkb4Z6CrN7X57TKfdDdG8hs
mQVUA9e7OdYfYu6YFq2D6VPJ6aMsrgPUYaO5gc4wk2POMOtYS/ZsGSn5/mOJoJ2pxxZlyMraVHZS
Hdisu8szsypA4q9sKpH7RLH6VptexzoxInpKN9KIpdD07ivbIPVRNTAkmm+qCR6zvyxNEzZLXcCg
+ThVxkbxEsFjhBFxVdT8nNUeB/h4jsqAznY1N9s/ZJycqZdwMr6S93Dij/ch4J5qMZnctIT3z0d4
J/Vo1ln9i7OhifbP6mWxDapT0eX/itXKh3b82BGPBdtVhkzHuzEK6S1/t74/C/QjPHS8u3ZFx2PV
KqE6o+FL0KL8QuU9Yhx0A/EjdK2yXS7X7ihm1sjDUkPN9NuHJCkpmJX1d1MwelPE2uwT43sVnKcV
CvZqZUrsuG9BmQCNEbDn/OR6N+xOSD3KhnXGamx9YHIoQhUFipaQNEPU55BlzKXMdyuwiPybW/E4
viQcSOr/YgeGOo7PKjJPUznUrwCyK4pKLqDG1xW7GWmyoh4N4FmaSF9BMCEIWZ7taIy1wMV+mbr0
HBMNUCCX43zMxPmpFaTkEXXYcp9XOty7E64DldntUQUJ3QPq3KlZJXOB1CTPDfOqGS9++FVAhDFk
p70+eEbkv0EYCEUg3+QT9fpZUQ40LE5HfwljycnQKBOWohB0DA7SphvHFUwu/9reZO2PCoUV6b2z
rBq6tAUFi40u6amWRJ7ihWIrpvWcwobVAu9SKHfI6NbXIwGmqCvKQiSo/PfSnIvjm7ZqZUvVOupY
ekXjxlhYWndXg6D98i1I5b5BcojEjEK1do3GYAInQdSnQOQKo/Gn8SKy6dWp1+/ecRKKgo1ywjsg
dh7036g9ZRUe8b0ANPG3+ZU+TGiG7G6zNmPQBXvhgRRxdmG8+kp/SesyJgoNul3mEUzP1kXt/TG0
oLDkWi3Xpv6UjSIJLBXEqylpfI2Okl1FgXWfyUq/WiMIG2KOGioqFqKB0JvRTcSGsFc40dSvvXua
YbvxGSXbrPhbMIHXrFFOW2LaTT4jEDJzuf5g6L6DjxGuCV5c6f4wyttaPu7tVd/Y5j4Hvg6b687G
mzdCzszNPWWpHFIReisu6fj6Dmkckr49qPy+7JoXj1BvKceBOpUge4GrE7gC2YKsUUetVwFHntFA
XRdhvotmydq081Z+SRkR+qkoEF6Xm4ewN2BcuUW3iOJDuqWReTe5EIqQYgH9ntyZ/mmSbP7qMqoI
EUp3jBHckFe7ano6EpiJkBoLQFRno1G9W2NhKnjBONEydmqGX4YiUIqhHku9kaysnwtC/lPdEkH2
kWcRBNvmjUuf4+y72SjyaRxzWAisEHD+3AzwD0Vq1nKWLhvPjqoUyYREIibVxdJ8dTer14mlklHY
Jia2tyFtFH7QDjTphP13wqae6yls2QbmGG6Y1uyWVJlG0LiRMs0ZHdWmtouQ4pVDPUoqka8q1PpT
vtEwxJHiJGPz6MCZBmfhjpFrYtkflXvvYMSATGi0T6IUaQgriuUM2aMaTBbwdH/Rw3D/ulYjnN+E
hGXE9gsobqLqVm8k4JpslAf7tRl0t5hArtkb8MBx4UmWj/0uVwSbcaHk1JlkZ3ZNXdaQ/2C5DCgc
NC6Aui61MLz/zUFWVNI0+L1/aNXZyYj6CwH+8p8sd3yPoyu1FlW/LX6B/7k/pLFWKSdOwcV3FTUO
EjDnyOyd70ATQyRgnZbNY+nC717cmFYwyiimhBg9nTVFr6YqSagPV7de4kTvlFwcIwCnQKdeuy+G
/KSk93WuStcjJS0TW+dznzDDVEZKC1ZP1ZhwrHJSgRb1tlV5NCIRQuxCq5kqwdQJFcTOrsBE214Z
IGzLD/yY58ALlVGdH2IbBW66TesmBC7IfJHpyrEdtADHp1DCRpTsfPiqp0bvmPwUkg+mynt438fM
/BiyhZFFsTUXqyxFypGpYC3fp41c/rf1l2yW+Im0yoKoMP4Dzi3lW6+92F79dU+weysTycBYUVq8
eRYvjLVYn1MIN7c7OsHusZTKUtzojWQLe/H7ayd/61rfwijbbk59GVnDBUrjoxFqUdo1WbK4oLaH
yzlH+VHAZ26AZl4DHaBgt89rRuVr6wZuT/KdBtoXqDNe4ezPERR9xHS52qoU8ye6/bp2l8IPsbY6
4+R5QKekER3wXCSFmwffeAFUaSedGNQfVMYiPVjtrbmFSEoLtlQ4t2WRnVvxaIfRj7qgF7r7u/iY
Xy4U6+0lq1LzMvoX/a/FF6C1MsFyQKakltL14N/RoV8ZSAwB5HiBu+cvU9aH6q7YQ1ZGsPQ9iMFU
9g2uy0uvQdP9znXGLrpeSt7OBkjpHuJeDgbDAKgZnqusIlI9PnryXJI4kUaw/g8xcBfA7mHUFG4s
fla9bKJh64jpvGdXS8sGWOrymoNhxvmyGGXIaCyH+y3QZ2Rswz198imo+VkbTxqhAI1lUzpBxwGM
NobF0kUfHj2Ejb+3lswmj/DgCWq4suTmmrT93mNwFhoq/6160cfVYRGkowr4TdNsGOUJ3lK+XkM4
z6VmmeWzSb6a/kfouxlvYsFFSTPWaA2ZfihvOyNCimCCzJLSYWn+oShWzT85eNVb0eDXSKta/TvY
xjl1C6iSgirdoXGLN7N4IQrv1RVvJrEpl5xvDUgLCcESDNShObv0igK8o01wiPvTL+XSrh9t5cIr
lPvn7ywDq6j6Bdn4OVTaeaVpj85kYv3O0nwcNF54aQwALjcePtp7VfgtF2bPqMUMt5AjYpHa9Imf
as7Q89peaCUxz3eN64Tg7rt+9Soo50JJKn7xXt8VUcxOF5VM8/nnMbVEe2dSWKu90gf0DT54iLip
FtR1Qe2VNvuWCRbMNp3T5vglqitusOpM7xBCleGXzulr4JBttqygJGy53d/OvPQaeO2eVjIg5ARj
O9VAFEobPQ9MZD7kqkvgtJtKpTj7iEtIIoavsbnyPOGLsMCndxFaUThm+oOM/orL6l75JP2RZprL
okivHsVCiWdHDeZML0sHyxs/Ml04iXIvVrJCj14krlsimKQeVsgXhKPxVk2zseLV/sUUYsnRKeYL
T2CUUwpPFZJ3v/BIoXCkSfX2zpZ/TXyHqKoIBmLbix6yXdtEINmnOyb3vNpmRrd3aS95g7WZiqVl
7/94irjvv5G+2trlBASdrWJ8LNV73i1rQYLPchLvF8xjgjSYZJYSBK0RY3UCdpnqZAENKWsFdRyA
bxvDnI3VTYxGzhlN+BmH4m4SNWG1kGCPdw7mGQePPk5wPMLTdzoH6ynFzcU3+NFit0vOhPMehw3r
8Jufu49xL/EdKgEtMRuMxMv2QlzH1VxlWvLe3ZW9VRLn9ALhCTtXS6NTdEz2UAAhOJGC6w5wvH/7
LDfUM+cNiMniDwstRuOAt7H9QUam3B4gICr8Yx3isc0adKbqmQQqOY3aH0hbrkuJI7tQS2n83DVM
NDHIRGUehxXOR0WqH04Nk0YEGKNprIDgg2DJmxv9onGGXSFsdD345qI0VIXIGqkC+F8+58ccI/+i
ep/mMLBBrVn3FEJE3O8yoKhQCjolPEhCD3+KRrATsFMpsiWEAVJf5lE+8fwriav48IJL7YeooMEp
+VH4sF9/VM16Xhfypt/RQ+Uuwl78X2GHXENNP92MdGGBme38KIg4iiwb7S3TJcVxm3e+g1Z83SLk
fmJaOMLKgaF76L9v1bKTTzzk1tlwNUmkN5FXfcBLfKvTve0urmwy1qQmHOQ7nWoWIOSi0u+6p3OR
KfzwGQPdDU/Qu7uJIk9wr0vFnduk2P67v17h+icU3h77UE3G9zucbsazTZWaS4pBVLpzIq/h+qXd
g9PAE8Yyjzf9iEXVjIgV3SkAnzdXDmMveM/Cv2FhOv86FVltD/cIE2E33uaDH8N2Yv5wsTQQ/C9k
/CsjAH88kKaXt/9NjeJKwjAOTjM+njPwk08KcI/MSEh2RwdKhfjMNJeU0JJ4TYG+Os7znro1FKKU
UHfq+PM85OA5hOkElWdciDDjYRuf5KHwm4tWi9G8mMl4sXcN0fP07W/4tNbjrKVcyGabHLvqUN6Q
gBP/fzdiNCD9b8GnFwrmnzsQ22jmuSjWKzOnXZwfDE6NGLSTUQpaV7vI0w2gIrmQJu7+GW8j8og+
crnUmcd9zBFSacJ1UWVH8bkJZaJeqvFFWqlV8re5G4+BLtIlt5EaQDgys/hZcfPRyYElgX51omK6
Y5TI9Zb/VS6rjBesfyoXiwIL1mnXSDF4BEUROwzTKx5MY8B6dC5YfBGoxFjbjTzNJWA3rY+u5fO0
CJn7Cdu6u0xMkmEDCM2kPFeOyRAUKZjz3fKnTkOiEUBbzfL5jHfB1LfC12Rl8zg8uQ0ZWEQpxBiU
rnWaLzirhxnAo0On3d45Dfybd3lkx2fMbJ8PntluNR79iW7WNmtwrQLT8BOIgUunFHmreRt2NQvw
Qus5NGn7oV8dyxl2G509CPwruk3O3094aeh12on0snJCqn4CTy1JEsR0oUjTCY82tqgW/jAlip8k
TDtmxekJz7iqdP3KFYXLBQjTx6Uvw4qbUqV7JgW0+zH1GzXRD1CyAgNstlCIvSun3G0suvFWxVRn
fpVWjsb7ZRezgv7IXKk/rHn8H/t5pNSzf1Fqh01N2ynyOE+pHgSidwsAAXsBmkvpi7iWP01ONsHw
AT6/u6Wp45kHwK9IsPrte6OG77yUwKR3dlpeuE0Qsk6qSnu4x/G47hldsIjA1uHsy3002Y80XJx5
lzi/47dFELdNJAaRPGIQkpFAfMPb2jp2D9rxwGTXXz86npItKZ5PDJx/wmOPJFiDJVDLutl8bfOr
0Fzbp1KT2st7r5eSk3x1qZ+FppziPQueKsWqz7Blp6v85mQqVVz5pKtdtW7Z/FVWgAVrslD7eSgA
eAXPNbw1AxONlYy9pDNKkllxPNIbc5Ukdh2/lqYIAN0mY4MD92eBn9GDoZB8E+SUT005knd2JY6P
LBeX4w8Mc7FzHn6se2rxIA9J2E2t6p7FQ3JBckxF1o4Dr4WewxQiSee/LkgXzsumkJXC8gptqTDJ
xNgwVFG3wgXrpov8z1gLh96c8/Jo21Sm2i2/pG75AUxJTFGKHZy0iQ+F4CjLdzgcpaKvb3FcPolA
JNiesqtSyJQfJavvDa37xFV8bDRrmsIp+cLep1yhyXBLTHEzFbBNwqoC7LVR8Rzt/hlp1JWYfb06
maNCyVD04WeyICslauFz/NRtP7ivWt4rune84hAknDZqJCbyQyzRE/srsVBLAPHK14CBY/PS+MxM
P8a26ZWgynpZmJ1cx2COh4uufI2SZfJ8XmWo4JbAfVIXDwGJign3iHcZoHivLPPtkSqFXc6htaIe
5NFjRO5OhnhvFWN05f9muuRoahbZKUNEBGbq4tIoOQlJCNffoaTdCCOtKdn0iXeLt1s1s9DSCKO/
vqBA69yDt5SAZL3BNQbAK7+o+LfP27uWnuVlPjbTLjD0yN3D6Uea2VejFlb9axZR6jOP5Do35HgP
3qa3iYQp2QBMJ6zLT3mhyCyeL8fQgn9Y2be45zJwJQ3YiPzOw4Aozj/FVgPpvWraz4ueBnPGCpYf
Z1IzzeD9tf8LyVppLhSkeNItvsFJBSDBZ2um7SFmelIJ++rrnaVD2Ir4Mcya9tnyHHcB+eZPqzqa
acpoP4/X43XJIMDT8E306aqtjSCceFTIdO1qw1h/NkGohNd9/jry56zomTMPjJ9z8thNjyJPBFyl
AI0yvYo4uU3EdBts/P4Ipd95Kx37csfP0h/EByueiR6ICmHIdTaopKm/Mixl8Kcb57LyxOXv8YjB
/ZQpk1T7l/f3JcpAE1SJtmHtCaMin2uJXehMGPhvTf9mafZiqJVYqTl17h2lwMrdS+APmoYfGHeE
CBYzf1s/nCvcGJ+TXUGeqzA+cYEN6tHlARHi23gcTgyYwjGrQFmnjyDIwnbqrLX54fLHIwXit3nm
cpimAKTE+kvXsRc/QztJ4hm1mZ42W91vrDBktrNgnwPpWPjf/l5cDOyyq4VtSZq2vi9sHvQhBT9+
KTBQ4z3DMSA7qJHjfVhr9+yEWlPO7xxhpIW3Hns2ldE0JfHGAYb72zUvsU94OQh3xIqjZy3lElCO
5IHHTRDn1fzFKEnF6msoMe+aR6j58+aFGyEg9xLkYBNcfIoR9skSsKBWn4HYiaiBKsnTZCdPddKg
Wjz1YcMbKaCu8NRe1OSVZDOQKMKeRyacdYcQItXRyI30qhnB/s5k/5PqrgOObKi6AvXKRfE/8i8E
9f7Luvp0ilB3PzZroWTZCTkV2CTAXw+OnkfVZk78oXDyEe1i7drM+LQ49roV3ydlxqXubO4IHO06
8GDmZIqUAYYBmOsfa+Mggsb3Mv43qHJ7pkSLGZwoL5Yvdtlk+oaf7NMmRRqbC9S0fBPesyuX2HXv
fogi7043LzpArf6s657G0z1z1YCJ2lwN1sWefXlk0UtxLMl5nwbFvBAJ90HyWIMJzSb4WwqkehSV
pqk1i0NdUfKGiQHSNMT/BKzU9URmjRgUIlcqt+VOLONVyRpU+Io4mGheVON0GmjM9uo7GZJOHE1p
ZmI0CmUGsdDSfNhmN2+dJVf55kDt7wJDjBIY5iaXnNuLxnjYuWbr6UMEmsj1TGboC19MCy9SN654
sVtY1DKZFJ+X4CujVTMTqWSwK6vEr/CEkuuFcIstwgUDKjw16liSwl2qz16vEboKMRQjY6Hw0Rxn
zyfIP4aR2iR0xiDGHefjwVpnAzP+WS9dLRnFnjwKBpZqEHIpxenEhilLrQQOHGoWv5/vPEOq+WMI
9AU2Sec+/rZ3os30yQ6vAjvBcriKKC4RLo2HftwaKmNXn1sxhU5TcQSlWNx+enU5mIECunQjXHED
NQbpgEYjbrEea2Fgo3R8yA7WxamiM/dMu88sI88AUM/+O1myyCdL6L42VeypxazVbsfrR9xkQct4
BitOb0R0pXzJlstLWuLsjsNh5BBsfgWNv/hVZrvDnuKtD4jUyvZqEpdwMBhH1XwMQVcrqGYHJ86n
MT5UVObFcOWSWjpbVbOx5rAY9cT/bZCT+ypd3AbDhpX7pf/hl0u9QBj+Ppbq01WbbpdtCZa3VdvK
7ZQcgdvwpoz1XfudSy9+QYRICS+22LGWujilPj52oerAZzdJcBa/QemFTH25156Fvl9VvXUxS1n3
fZ6dAX+G73wFx0WdyThXc2IHc9wOy3kLlvzsxIj2Sk/BArvr2fxKtE/EWdb85/JF1x1CGFxxYgP/
Oxvc9KbrjI67Z8j+h5OTeAOqhyazcNjvLq76M5kIjFRG2XI4oRzP/OyyqYl0gOSwfA0jvBU6zJNX
mqfbJsA0aJmDseUHKugXEGTnAkejm/ZwVck0gU9oyu6bjFV2ZQ92C46FkiLxYpp2yeCcukdTJ2g8
hyLXW1Qo/vv3NRuAfUAtHZ5XSV4c2NJjhJDyIOtAVe33agit/9vX0bqD+PPpiZSxOzVKR0imW1Xt
66TCCVglsLrTsf7w1EssSOIFW/PpfsvbmhqVgasam5UkruZBiVG/ZsBm0vco7xskiKJmhlTIMu0b
+ly/1vd+LWlUThq8/3ILORcwb+Ptttc86o6J4FGH2J+a+Hkp47W9NoL4lA3M7B0loCE1QbMDBLIL
CR1SVzxgm8gvEinZ5QF4+cx2OT8M66d0hHf2BDzCnZHqd05ghUpzsvhXJ0FkpHS2EjdiqTFcfU3C
GAqjCCIr8WN7OLzYnS3xX8NcjwKTBuTf25hcZJH+1s4YldY0ABnkbZqwg9LT2QHlLWgRpJPVwjrD
hB3/LcN/Jzc050QnpvXLfNLIC51OphFl9Ec21WodRK8GXXP3lfqVOTeYpAPvW2DBibRkDGBTIpPW
jhG/hJ36b++xKnJL3WN+p7lvYIPBt+dX671zzgg97LRhfpBh2Y9jBPjXEv/L1Z0hJjhewmDp++1W
O3/7yjLrahZkhzGFTIwxXaxNT95ohHLCXG68h4raZeUa6pk6s38hofjhZQHMfKEljwXw5ru6Rfew
Rp6WHDB1xfenDPflCgtuywtPe1rEt5mfnmmDU0rFkpwTTIuxYIOwUnxKIFCciWx2aiJmRtLiiZfN
vjDnckU1GJs3h4baYHUkjW0dXvKMfoPfkZDh6muJ8q2HnHVbl7fGYz4zCogT2YnfM9cYcipcvs2D
wTXQxYJ+4MUkPimyoIoOce/RDrhAMyv/FmLtWlVkRKIZtBZ+102I2G4ubFb8O5mx35TAsHBEvGHL
DNeO/40mBm0PmbyAr76rXm/wLcp2O4OwMttMmTFtzZFd+hjKjs3z/swCcbYZz9gVq8S/wxhJlf0Q
0YyJPzEFDzDr5WCrMfPaCYLs3yOnYuTnDVfsRxQ7n5qP79Rn6IzxlGRzZcGl0HJKiwVILt1Wxo/q
v6ZWS8ghoDILS1N8aZ84Qt+bPMuf9mNWzIEYArPqovB0E/aBBHLtE8cWfCsWUHTIp00VAcgDT8S2
DwkjU/p7FA3IslkfH9l7MokMmNIVVpNYG9i/QArhHX3sBIqjF6fGC6UR9azuWErd33AIybkV/jZq
WxTeduu1M/nTxBsBARQj+V2eY7pWPbfyk7coTWBx3T2qau8KtOGiSKA3Th5Tn9VBopymXw9bFKFu
M9qvMFrqriTdPBEwIgYj8jIs5yYvAf+UtH5eQTqkHn5YQfRV6QqJAQ7OS5gsItccAfcA+s0Pzssa
T0O7kyrdM92YYwPyn/9soJ37XN8xhqk366gi0Fq/EvXIwME4dhCogUkVe16/YPfg3R96u6iZUFVA
blBa1ZtQl5ajG9YVqcTv2w+JT5vmWQPM8Q7s8G9J41M+qUlvztcQd19mADv8o7Hn3JoV5hqbjQAe
6Va4uJfrktqUzKu6Q3DCxBVH5CjGsCetyu8Ue4fGOX9N1Isx9icJ8XTD6hePuALvc/xlvbd7hKg7
Eg7wcHrp89K9CgqzsQh4oeP+zi68tfsXx3PbHrQNi5EpMx4AZhWp18spsd3jEioC0oKVZk7Onua4
+qnq5gieA7GbF9Vbf/7D5kkuqq4+EYrW7ynUA/tFTJznq7Pjx7R5ITo/vFaYf7CxQEnpsmyGY4cB
I3tcmRvRhoIDGxcHmuplEapWa0oo5kHWX6msnfMlkIuh6hr9FjbE+puLvUEmnmssVswKNWmmPE98
bNaKo07OMfutGBTtkqad6SNPS0dcyJQMDaUkTFitryXz4xll9qHxPkUkP1JYGjf6Tn9C3pb55CmK
5MkcFigJzEPpZCOOdyhjpCN5jHBQeqzJKWHeu31TTMzEYnu2aYF6Rj1EDlmCZWxQ1zzYczrckd6C
8b2luJxj1PI9i15fD/z/+qW83bIzWLDx0MBJv+WOTfzJ0ajTs2bCRtKuChGgxvwzK1JZB6nNwVHn
VPmoswlz9FJALIVNjBqPWARCHlK+7KCPb9a5OACRGXhwjLfNBb6rVaWx1rZE6SCEUfH/d1BdUFEJ
xOJQljh+ik/+WG9P3rGCID1WppiOZa8s42nq0ecM2hU5GFbaq10aOLFEgzqMJzBEPBksuajxWUpQ
0p4v+R42AoHNINsCa9ylqHUDxk3EkwZZV3u8yqVUir6lX5YHc+3vIpJaO60k8IBTL5oH6sFlVHVd
Ol3mfSV0T3VrHgQ4CSsUhtPOgHidBXB6tqEIDmupf8n/p8t8fBl7XSMEIikoQPbio0NF/72+pn/Z
Ek81ZZzi99dyHDQtDbWe7YgkYi/tZhia6jB11AyjOWEqUbpqjNLfkgx6rVdJg28aCd8wPiZT4Wh2
/8giVKh2CRPgj43ExgEBzGDRImySGFh6qRbWVHJq9At8WPQFySA6luTtCdB70ty6eP0dnXXmEenM
tNxqDhWa0R83Z8/qPp6gVJNqz1HseSbH/Nb8+BfJMauhB8FNv4GCMFE/x4WG3HyZMDnre0tsYnnY
V2SmCFfn3rn3j5LeR6wycdZhtoSI1vASgb6/z4FiGhaFYiA2qatUHzLrWZEZKH/onV0IlgkrqVrc
GY1frCeu4Nn82BmvdHEpGTYnk6zYeM5cpsG3aEmR6LuGk7yIRclVSNVuAggO6zpFTJqN+vztXEoU
SA1JFgm67qSxc5xwoDy8nFOlBe/kJGPn2TS5soD9FkjiGv59kpm38bcfIESGYeC5c36AK9YrwcVt
vVwm6PWBODbrize5oFRPFPKX4EuXuV0qllZ7XwJED5KqwMKDgwQWAzPKyESqzzpW+XxtNP0mCoDT
huGZydMUIHsNM35R0W408cd/pyYU3hy1cbgUmnv1ILGqo+d73iqm/hm1Gn34cOBPARHcd0RUv2K6
2yCLD8cS/HnMV5ye1mmuvAkBWPF5IXCbqO8uNx7qxPDeScM7WKd/2CPTIanz1yNmyyW9B/SRYLXy
S7TkdvBLUHnfyLZ5VathHc9BW+BS2SgY4pwZf+dXEGoaM0Lp5Wtyu34xkqMjdXkC0pCL8BuQIMEc
VgmiUJRmBX0Vzxq/YFitfHAa2BgN7Wbm9eihmFzcWck48evXuQ41X/6CPaaPzCorypbRnURr5rMG
MBlpO0c3KL1zDibKDGDAK+jnAdEAXctrbhcjeUS6wWZvIRi4upaJBH+A6koXUn2wbpnbBZGZ6LkB
3FFTLjWIUiIjnANvL6IXcd1IdvPBOxjqHZQhzLaErj6nbYDdIkp8kfg4qwnjIcXJO8vvS5N751il
tY4ODfVK9Q6m9n/hJIKvJB4qo/RH8gWXZP3FrEMVgf9ZFS8ACMvNl25oJoc4XsJlF6jgbxpIiIC+
jW9NHH/ilgZ6phSA0jTBtk9TZcybBX30jDrlCe6HXM1JBTpPT+J80CFHTfgumQhmMw33A2gzn4RJ
8iM99mNlx/+VR0pc25CK8Q/p0h/TL8+vhWylcRs8NapzIAUdYNw6pcL2ZI0bCQI4OsK6pJBQrinR
OZBy1zPxmilb00jKfGOhPQjNOXYPJ0BZdiJz46zhCf0j8RlIsieXSh3jIAxJi/UxvMKEyL/5N+O1
RwaOGTXPW4VpgODR0SKotzLz7OWtddq9M1PPmyzvzLeBZ3v6u7INnKEILSfFN55yLSUBJZM+VBxm
MsM/+8fSxsbbXEbTSKOSoXJbmCxM/kKz+ThNxl0TapPbXTKlElXuWjjnG3Jo0IPL3aZycMmwY5Pq
+pIehwcIT6scdBRkMnTIegj5MM+cuF+HXmz9fW0KTjaFA9ORy35NSepZ0FOx84awctUkxNRtqzce
leAx57ybFImDLjZVEaPF8kIS16XDFOpIRs7FFBQpgyGqI4Bf1kqtRCj/pSGsFFCDpa/fZh32aHRi
gBVExSf8PZajXY5fLXZ6Zd4JweEY4ay4hCyjamfyncrvzoM2AUthxoqBmn/r2Rd3LuJJeBaLs4CS
ALbS2verbypsY/pML/HEMqTn5/KzvC95hTcFFfMCitt4JdULxfD3oIjuXte8YcauaOvTTSRyhMsn
lYedfjVHQhxGESZoKGjxPN9UZoAn14KIxS3pdEF5RTn2hzEmV4XVF6vnGFSK0n8YQTGent8oHduO
dqvXA+21tg0R+nj0NBvrXh4WOyRF//I4iGtrCxjSOW+5EIwVnB8j0BmZ98iP/LrQJLOxOgSvSpzT
z3IWHXLch8eR+duaT2Khj1kvQjmYzkYRSuhXaz1f1r12xkdaJVb0vMNNOP+sQ0mzFAaeoXhoECMf
t25P6SBl7vYGEs1HnwdPdODfO6CYELtL1bGcfBgBYlzMsyeLn6dixQYrmUovt1LPYtuQYvcUM6jh
b8SJREl9EK7rHiKPRvVBrXSg1xY3a9DT2iESr59EiYjcvc2WDaZ37g6hPDXF+jGcp59Z/JUvhH7P
U06OuPXbqHK0nR3oWNaF3P2N6vsEtF/kE8YWpkljwqT6Evo9pe2o1vl3h9U+HxouPF8qCZ0yv7IB
fVZXD8Xl30DNtveXpsY6nd00+XXrnWifn5xGXZ8PyB71JiUY5dKrQzGeFc33zJzoKKwARzIu4D4i
M7KLH8jA3zvM3pAa2piHlmtbibPBie64oZQyVvsvoBQvEXUTaa3GhNIUPmu1dmd7CcErmS6q1V6Z
8d73zgYLXUN+u0miiqw6XBgoAWw4u1Xb3931plgg6bZrF+z4ose5xPD5JBxJYrvwf038GVRkPL90
iT5rFqGJSosruO15j9jii7tn0u7GGkGZ/OvWdQ+quARfZ1ZzMSnhdISh616OnVdWotJhDKrzy04N
Jw9bToYBWIAtHTtphn1iue5DU5odLskCAFRe7fY7EfATV8mpv/Ts+hI2nNwB574iMDChd5MjCHZ9
0yUjyOxxeEvKibuGls2aKzpHep8O2e/VIC0k2PvTtvSTIKNjv778RKhwlJPbVoGESKavIDE32IRg
YTTCiGwS8F24BrVPhGS4A1TfX27sch6dZ4peltvMgwNwb11tARIjy7EKBWhKxKdiyK36on1cSVTO
jgSLAG1X2cycafv0NZ9neE5WH8D6c+vKoss1+9KugkrroRF9HtEKyJLFSsYFRe/dAmKgNR616Ecy
zbV2yEkUmSvxDmvyztaBcaXvhLxPRjDqMSQPIb2WzfnbXC/b0YBtaCzm0C3nINmlgGjOwJMjk4gw
C+z0eCSt00aaDzRJdHCUEghsjQN/uE96VY1HTU/qL/8QNc5MydJNRWo6HRHKTlTbLkiiKfPlUqk1
16RuEQC4ivn2u2ORHVF66tselF2wMa8ho/5Jy++mdVHtEsrn85Yklom5xN0uyvP3OFGD2UK52y16
sYbVuHWC4fASO05DT70oJU6nxsR1mtiOen7mTPdWNuKNUYTBZQCFZheUhqJj1VtfXKc4/RDqzFi9
zpkvXwdLhOZCjsyhTF8hcYG6hIjPTZDpfnJV0JfMPSmBRNBtAdaq/YWXHz230Co1DrU8KQ9l4Tj4
YpBtM7Cp+1UmKa8YO3clutI/7gHlQX2Hf2HaLtZBv3PF7zwaJZCsWvoWZ/ZibZyESvCk1/aJEr/n
EBsCb7V7aEzooND/Zg195HPE+q/pJecWWLg9jo8/il184a2epnIki2vPLr59o0ZvLgQIze2obY3c
t9VLxXg9cX50qqDg1+tjc6OBbahVdzZYwE2FPjPr8z2cJmqSySB4Y/hshjRjPzZK/pLUUhSHUi4y
TKm1n9T5hxKL4GOHKxr3vtjR+asPh5BykewMyT1bHkyyY6TwfdsAohRanz2bkKWIX07gCGvkOI9A
ahXJTUXGYWa4eL0VMD9bWij207OSaQBNIeHo22piD1SWxix4O4gW49a79TMPaS1+alTbea+4buQg
CKDmuCSLawKS9heq05KMP7yUVlnu9oSUu/aYGo5jABeBY4vktkm+mzNRToLdHQS4My1y1CWbeyR4
3WoNEAvglF0hv23r8OurGWCJoKIzUMrJSeb3pQEeerQeyC1j9UlmJKAJ3aPB19WgvLsOcS1526x6
9FVoFYaGPH2Qlinvm4aO3c1zK1cSXeNCe2N64XvsE1DJ0dc+v1+PuNjqSHUr2YAr3kqmCYnAtGb6
wSYStkIh20g7jl6DWSDkcOiumkOEVWYN3o8H2L5XWRo+8LWolJCYOqfxHsoLAOPtDGoaeJZgHpXV
yvVTNM9ZAvVO8714TMf1WUxjwYQsyPzxJJ1H6/zfiC40TMG0fhyAjU2PHTJyvAzZmq8WHfGBaVqr
9HF3k6ORz/crBEFt6HimJVV0mdxGbrl7Bn3oxOukHl5HA2mID3m/46gr95Oje90J8fGwbXz0jmy6
lt5f2X0p7suhaL6Y36NW32DrMSgypoWNYUjBnHH+H1JpYETjGcamk8nNMy+XOdSLXV4X7n1PtwmO
1/TRwXm1ht/ccY2eyJnevEJcSnqBi01f710Sm1WRmFXe6y533mYZfuB+YQxnIOnrr1sF7yn55nyp
3gjQmZdiNVeYCTBoXMzYiPFchgQzzdI/dmeAfXAwjfKCKqHMRGgDSD/Lyb49n4LkQOIPKsWrNvB5
jF8ZhL9+MIkGhqBO8yfz40dQME8okO8fCgHbu1GhzbeXhtW32Dc+gRz8n2w0wceWQ0ubRGG06JLU
gSWmB7JNS/da97s8rd61FIsahgP9A89S5eRVk6sk3vFYHLAmuaxbLNpmkRqGBm0hdWvjEl59gnzF
8kLOvLGNNX+1rPIqRoninCVaA8OGh/Fwkq2KtBnbeIsK2LcrVSi5RXiPm+AIwEIGbQZQGY4VrVFF
NTgu6SnmNpfRseYu3T6h2atBZShSINIHebfKQAR9lyHqdQMNfh9z0xbaq5doZ54mccvJDfDq4zYz
mwke8f9NNxGUVPC6mJTNk0YA3ywq1SW/exzcGEMzgU4LVc+odl1cc3Yf0KD+aB0GMqlCY5a5grZm
DVOloSKge+Mwpzt/uBFvObAcIn86WOvOnbrFuUrXA2Oo52roXIsU9PtlYTcX89gGbMpl/tnSzKz5
nel6JGhODE3JtrUnHlw2xIbnd6SjGWydCIgoDtBLKNQDgWuT4SfVer0rdwMIRvd7paLjOFCv2iIi
qFC5i35K+f26d2TSxBQOHn9GLXyl+/JEMIIAGfIKG40h3+GQAzsiXFohMi07cvA9hogfa0nuRK1F
+a1HoX1KoEdY2G/8+8iTzX2wt32o1G4rPReQ8uDfyTuQ58XUcGO6YGY36sPCprQKhsWBi6Jqgf3X
nrZsbCiTsk9P4l7Zu5oDLQPWsLtjnMHCe9GY3hab+/zdzT2Ht5nHXz2oZnolZhKLHylFzuNv9hi6
lV6HZmh2NN9TGEqWjtVBo+lu8Jce4vq/ZAhtZkuGqYiducXsDMnhkT4xp2w38TciwWBUBridVf/E
u7p9wnDDhT31LIXgrzIBUrrqQxJRvy+nxSiJ/8BW3HWCJ+c+vHHF0KVAWitvThwDMzbiOXfJj/mf
QQJe6Y/Hd53TWRGgUEAmh8ffroVBt2lr9ZCgolYsmZ6hL7zwPxFij2+Hig/feq/Y/3yfjf2hWvQN
SrBRgK6ymJAJ7MIo+DTztZVSKzfWGedy+DVy8OpbJO9IfFXiO7ODAhRYWMSPBsGqux7JlHwaQpdt
GOOi3tC1SbbFRZ/jGgVIp3b2erfZa1hapKmwFm2IeWDPraqyhQ468H12hqmeXoqOfceARb2iYPzh
90dic5p+5Em0r9cKi9wia9JZ36rc3FxDF/7Mn7oLXuB2EzzDtKC6QjQxtFkNVOl1jGINyztfs9Y5
ow9jYt21/1buigNuw2Q7eP55syer8GVhCeDeoPuXn1zXk4h9ofuLbH7ovsVyWSdje1+m8BzL284S
QSpnpgL6NsstkoNljuNkd7OfNumSeFG2AXNlIKErvn9FjDiu+tE63HWfO+dg7chLdxJAuykbVecR
Xh/ub7kZ9y8GwJAIHmUL5qePOGWCsqKGoY07tp/uKob30EqpTJ0WBcLWVvkuWpBkqsexo1cvX6px
hYQk8CT58ys2LUqfFMikc/FZk6qT7IpdZcDUFGRVPRQMWyJwT0MZuuz2JtjBmvY8vLGfKPsvs4Jb
Hqexc4FcDM7cyKClmchDJC6QU6j0chxPxf4MJ6i44bhbe+yCV8vSCRev2/gM+8wqfLrXe2dw/nIT
/Vg9RfjQ3UYndLxNuKfJgRXRheAxCkj5eKJwMfP6hwjTkkEnPRYsRFAjkDyIRpjsFcgWMGwhoNsj
HxksKXro/ySp3itHoCHZqoqLDFvXWUMJyuOaN0lh7hkxTP81hHFi3vI0Hv9P5CHcFowRnOXhNNuQ
pwIpFvs3niiYjhVCTf++O3zsbEfKZL9AtN4merex6nqQfSC2FBAtfqeeAKYq6cZLDbXOZ/9lL4qa
MbmUw8rPh4UXkwB7Sx/ILUdsWQ8iLq1TcSsYzrxu2tLsDQhd17X4BfH2awVnQ/orKy9nLRHfuSvy
qfhvYA0ki6rmqdYrNM3KnlJ+M1QDdosyW6kFQuUaMt3oozrsFRvTba3mTJ6CZ3aHs7W1cQuozhkx
LScu07q2c8FR/19dnGXXNHvbsJtRYPdBPqvg3Q//sUJnTIISKl9ChZ+L/Ov7A6PKy8p3mMSAlY5v
Sg6cJKoSMAU2STAw275+1izuZdbnlz1ZiOx2oNT7jBdXNbGHgyPKUTIOIJx8lD2s9K2pZVmpQSDO
rfTwvIh2RFvHQXl/cvTXZZhaCXlSU3cuXNTgUaH8MJZsFlMROH1ZihdPJpPxqauxz17+8yvpGhb5
0kOkFKD5jqGffxhKjNmEJc60rKPNOqkpIvilJqQrOhb3NuyGDYm5Cv9KHc2rdikLgIYjcx7Kr+Q6
nroiekmSDXU/vKKPAgj9oRiJMdWO99wgKkQcb7yxA9143mM+NIHBXyQvZliAfRruk+e62i3PytRQ
cSOQ1GKRmDykD54GpjINOMuNjPjg+Jc3NcbC6iLh85ZHAbGdiivC/DfdYqcPl5zL7WfsqWIpiSLj
uW0TJXL9lJytHmv22WPDsSo9DDYQYiSDSdNHhQaHuU+yi/FfBMrw9m55kkqKxCLGE5Tdqg2s8v19
wBjCc/e/iTIBkeMBS++5JFl8Mgext1TAj4+0UbpiuFhY/HX1mdVJAR64FZG+3t1plc0X88yFWo33
C7nDFW0nMLrXGRFuXCZlflQNPl2+kAXbAKiAanSZEXwqqah6miLUZLRVp89dtDudhANDk6RPjsG/
4MDHtts+wQlYg4I0STTx2Me1Tqa2TP45f4hlXQ9ubIRFn9mKlGaGis5iMDVVllh04U6S8DaYxAI4
32eY7raqMUUFQjeqqw7j0PWrSvYaen82s5t+0K3D306iE0eI4iHHtnsLEMpttPpkyAobvurn3NF0
c6bc5pBkaOAMtV8x72zL6zEvZjRSv6onguvGlSlzR1X6tY1ON8lrTNCu5eYqNLEWxqP5E+rf5H2u
MTGJnF57kmtHIkxJj4R6w+pTaqffLJc9k3imfFlhIS70Bjl3oXEpa5fTiP0L7YB1Dq9yTWYzlqVg
EmrW+wNP5n33s+a1QBDVSTMUhkxEpqjOcvIrIzGrMAVuvX12g2p2B3QX8hn/z37aQCTt2DLpmp/+
27nqutGm3hDGqfyJO46Y4rDk1+p9O9laAqbYvk6lsInNRz4YbGx2Rs/KynBm8JGRuQjtJ9cuSuq2
gmQpSyTFzKXeZX8fI/X0gLFCAAfyQt/zwo3KSOo6c9Ejng07yFnrMBrEHMUDA7N2WtrlmtOSES7P
4ZGipJm4VkG4NuWBEtgx8oBzE5VrJj4AOyxi0ovgqcqVWqwTvsMB2Kdev9tQ42lJAQoY00l/+cdJ
QeuQkquwPBQTuoamHwpxHuT1eu+JXIKjcSSXaZmYFYk/Ao9BAi3017iH+gfiAaAQIYKwI1ycO/qJ
fFppxs+k3IoidLzP0Bz/q/zoKpOHQNsypQKuQaUxR7gQ7vgFpkMu/Kv1iT3HN9YKrc4mGJ83UFyh
9RpTn7dI0rzw6fO+xC66l/GnSIMKng6NHIpUCPTSLzXSa5xM9XKK8MV7X7oOoUt3NbeHITb+Cj6q
urYd0MZuNQzN9sxb16aRGJ1NkUBGYqd69BlO6K0QrRcTa/6KxAylsJ0atAkrKMtWMn95ndKMAGFr
T5Fb1X0EpxFbDshWghmcSyVMxzpZMtHktXIQmMyV1glOGJmg8kKZN6o2LKZ7DelrDfv3b6m/3XoA
Gjj+1suKUbaR+/htx25dNNb6h5oOjf1v/jiJU7Cu/o4STKEoBjIPoT6EjGForCvWNxWBCNWl7D7a
1kvOUkLPNI3+R3C8gY7UgO3SjxaWP0JraeXun9WdimNwC1NuKlPmch3VIKG/63gDJPhyL0PSKvki
OoUErWTXT9LcZsUYUaM3G2U7wuZji+y4d3jVo2XnJCSN+tEIptaimhvjhcw49bPuP3VwSxU3qdkB
7B8FmVTWN2ism/8CUcIVt1WOiUQ2m/VLKm6hkpEl4mKjIsByPlitxqYBxy8Lq9DVXlteWlaW6z3Z
oJjQYUt63nidov4kzt/zee7g+MHYkSqR2+98iqw9SlTeJMGp+h08KTcYoTHBZuRP2CaPENJYMpms
rl4GQWiI3/k5sxgIhyjKrPz27iDHNb23XgZA+Wt7hkz9mSRg13YNc72wyAmskdUtmGD/XJsALtFT
qTL8nO9oqOCAi96dFYrlpoikuXfrO5dDgx0Zh02DSdMb7OyCGzb65VaPtp0fHSRQJS7fm1Gugyzd
VTaVRWqU5vydYQnawoF4t7/+sghgud6bgrlTaIPtR5+1aFX6CRyFkChO69Uml985uSbh/Dulbk1+
L/EUNI1c93tb8XWQLVHzRd291iazs8y/BuqmmSHj/swMPu2FnAI0N5TBMIpZkOuSSTOP7xjK4RfK
sW8AY+WDiH3UuAK23MQQfYB6TsWzpUm82jj+sCLjh3F1JVceA4i6VecD+z3CNJd3gXGTVVEt41cP
NxFV611nMozasjCQk8NAPrSNFthJWOjNxdvqpTP1CaWN+iqPkAoSGcOP2P4Mt2DZ3SEdHfK2XN7Y
QXiXlT+y9o+6EpKNJ5DFj3Co6jBj0tp8vSFKJklL1FLOMfOcXKcJUKKm9t6kkMXHBgl9ll6K5U3I
ygQgOezOnSUacGdok51aare3XDPSZwPoQdTCcWuRcdkx2M71sNYz6C9usFj3J874t6HuKqrQYAo6
QPEQYXmk9XJCkp/V5EVMxEjMIPLeH3Mihi8HfJOherZRqRlSxldYhZiVIWjWHLwK9N6ma5KP3v9U
85vIuB5kW5eJLENLdr5iO93DiAyHVfs6IUOi+OHO1JBVHqX8dHmjzRnBb2IECGjrMFRa6NAav2/S
blzjuI+tYI445BKdDuUJNpMkaZltRO0tfwPT2wkYOetpinsJAnGOOMavcY2wKNxUXdQUXt1v67ET
IPN40hqS4qZFdMnPpeopdXRNslu/m3Ob+snr+VN7VEaCnioQaebhs0RFrcima18cScoAgOq+ofsX
MOQNZHsGD7990S1nbW86qLGF5ZvEiMPpxCe5tyM2bvyHy65FbwGZCZ/p8HAgbu6mmHtpo/fcVbUX
ALimY5L5J5rbM7mQZyqpUTVSiy2n0nYrCl2i8ZrfiPGWo6vw40BvwTn9s/R1eJL8qxaikO/NylH5
rroazAnJsbCU1Axhf33UzhH5enG6fUA8wleqbAWoyagnzHgwKPdP9fRO3unFNiMG+tq3ExjzPacr
s1rCyN/giC01aSah1WSp5D+Ux+xXYAX8Wl4HNeoEvlP6qjH86aDrWwLaEgMjc71aoWtrC2E2RPZu
D4vqbl8x8eWL6AlsNoGnen0tXf+sOgrpPwRy4zcpTqV9qzvAniP4M+VsThgHPXdQzDbPVHs1ibK/
YugHYthfMUn2JJd1E8xEXvfyFyUbQL1vd5n4lxdwyDQAW4V4PTQBB9oP1MX3PYq+Xx4VbwS65xEQ
oeICEQfy1tpmAEwrmJbWvy5OXGD8Pcxbmp1vD902+bwR/W/c/4FWkvNWqNgy6LiVWwxhvjwqAJuV
Sxf+ANzTQoGB2wu0P8Q6Gti1Dq1kY+SZsFqelrrsR5cNLpIEKDZc5O0z1RsIBM4F/92HHQQjGR/N
/CikHsNGGFKYJkTSRe/GTVbzNfW0gIV1hJ830Sf4wj807g0NVshQkai780Vo/zFeDHY4TmkVwjTs
a5AmMdv6vrWtcRqNOW3CJ1dlrLfcyDyFOpuC6/yfRqENVy5US/m3DXC/1FJkBjsAFWrs6oqFxd0+
U1kljlXq4DbA2TqsjrdaVIPp3flg7qmjNRp3MX8WuESKucD2ofnRRwRJ2KnVCBbaa8aYDcWH+Dyf
yj9fxi9RHmMAM++2z9Zf56f6Pi+0LYAXuHbPS/iBcaeMF4iNV8t/3hj1pNK2Px6uGd8pxKS318Fq
plHvLrWlFy14xSG6aSGC1MQdMcEILXq6Yn1bpGSKbSvtKPNJUfiSisxmIBUfNf15bMutLGoKHh23
9JVBNwhUPYHGX9rgf9dboNssQddKx/OlpNtnnPusoVUpnQ4v5+TXUYyyzj5l64u8Sz07/zEb8hby
HtjhD9ogv+64610enZeO3vvHbrW5r35yvNTJFxOlhlYMhe6Rhcp8iFt/MZd1nR54b3wFXoIwTxbB
rNG0P2nGdU1BCq/lMi1Rb1N/K7nWOGvt4006OiKt0CbnFGpRQ1rwa86ZH3rF7i3b9Pl4FJzeFj6O
VH9Vjhksngz67JPVB9/a9SxbkYTyjcvmwRbP4EofgmB26RLgXUP4xbpr9YyMI2RbUwc/S4RS97of
Gbnx34wa1lbqWCgxDYLj9w797EX00PQM5pyXeYkCdYFplaILVNj2l8PyRkwTuCTf74yYrnx0RmPq
yfgl+kTd6G3iIaON5WF/3CD1RMRUimg9YWwwNnVT/DFKFx7WDi+fpcG3IXSZhgvAOuEKuxp11/cx
V8bXl5sglavC0bYEyFO9rZuSqbMjoKhBjWkr9H7vvwoxg7ckvQuuef4Y30XALmTKKbX88CN2IEFV
v+XJyFpCW+7gkXpz3OcdJw1CGox63+INfNZ2UXIsKEAAbYwg18EG6aAc9rQcH/+mDw167jAcpB0w
qGllTLnYIxhz/pG1sstNjBhktOEysoiIkh06wP/ubUes6DbXGiU/04bZArDx9bIzFSDJM2qdIKoN
xDdd3gbTS15RTeDg0SsHlSVvd+Shu7/7oOZIudKax6FRWglg0uIruGAbaNZy/ZSLRwpAjc0s1CnG
WAOq7fqEtQgWIGDjGzQ2UVeax9tkKj4WTNaG9GQ1N7iHeygmhE1t+awUdpuaIlh7Gn49GKUBCh7V
JX1/X6J0CWp0XcMw0HR7PuYd357g3gfZejkDrXs6/CyVv52RbQlKzABFwsY20c89aBY4BDdoGSrf
eSyWPAozA/r1eBoAcDilVdVY+3LBK9kOhcNMuo+CkAnGE/waHx3C2Gy0CyCvabD9pGznSJjkjQ6M
dsrvp+TKEG+3cWz3QqTS4NnVQj1l92pR44KaaABYqpj9bOKIVSEVTNfrmWy0RddVqxTt3FmOr5Y6
T9ymlfqiNmW6BimMGUQwbt1Ol0aKrI1b5pBPpLFf56tioKwX5SXYKkrLa2Xm9H8yHLPbVbAB0Jdd
3eZXC41isKOABoR9hlE7svr9exChp915OJzvHXGB5cgfK5Tc7ih57ZmG3RAgu3B3BPWmuZHbyrhf
MzjZhuiBVZNRKrKpuCixXCJz1aRI6pOFijISyCWoKGAAExjixoTgE7rLBx0D5DqlkAGBvVuVfbmr
ebjItQA2mG/UV1c8NAMbVf3VJ9AFjjxJ6/AAHKA4ieUd64kXm4y3NCjO95x3E5iKa/aYucvYENwQ
5c044tmhoMNMqvx2Cy1A7be4pvCLjSnj74guojnh21MZp15F2H+Lj1M3D/DQ8JCylzJ1BKFp8wbV
uXo1rvfJRvnaWgzXXthUcVh8xizgwfBnn9jF8G7m3B40qdUEUL/9XV29q3pdHbAO1NZQi/4t5l3n
Q3O0tl//49wr4XIIGdNfEWaMmxkxK0D8O0sEsEkOKwYbNIRjjWIaDfnENMn+ICzuvnvo222cg+BS
x/excM0FmJW3ckQh4TK7oifi2uVEBIZlbfLRZ5dS2BWrbmkhrYrtDKMjj+w4Q9OqvBOKpliDqjzH
b4dVuvnNNssMhVJ40v8X3GS1+g15+y9ifFivkDstISu0QLV7l7JcNYuxA11qNB3GypKPfwgJN/DH
wXg9HqGi8SPWlI/PaSz4KK/YtXfUyX/fYpr1Kok8+yJPmwsktQGc01wcJEfnu23rJRZPuWQ9iubf
+EhH684Uyz53FVXZT9L2wAYwsX/9g1rKn2xLvDjLKv89KCyGcTyP4EIwFXyH1r/0yrPgk3wu5h86
4x3b79mMjTiQga8UCQTcsKxw4BAVd5zCN3hKUECZLWRtx3+OjE7VbPgfKb6j1aqPo1qOfdDq/4OG
a6FgvrYVzVwHQdthVQD7DkQbnPJ7qOmzqFEtnPpZKP5NujyESdDtj+VYTyO3d3Ri9ak56yhE2oLl
b+mAS4D2G9e4GJxP1fhCE9VOXTxWOB5acbA5gxdI7CUIMC4huCYdHyA7pRzbkSCrCR28QMO8MWCq
BEUhV2EUQW99Vc4FclEhp4eAFqgJ1Pm2mVpFXtWRWckgrkbAR3YmdQqF4ifGs7cHrZgbFsnGb9Bp
ozrSYnOmwQNAYfeuGoo+PHGSydr7DOXSJExUvygrbBEHL9Oes9wyyEP/qiTojdgix2Zovx9S+KLb
tgm60rV9DeLSu6nefxXjQjpYFbqE9Fbjnf/yq6SZkFCHdSFa4Myn5SpfmAVk0nliUyanioJUZRv4
2+SrQDc+bQA+9cVgakoQzSzcXco5gVv6WzkpQKGiWhmXJec0+Za1Lyr5CBdEZWR8NMyfP18ll02T
1+BXTeW4b6yuLnPW0wDrzAcF6ZB7HW+2oaiATTcDcjs/uxVvNKdsNpFTfYIig87ESsLD2MzVfClx
ug8jTO2PR06xAsfXwxA/ddNg2idmC1P2syXqH9NGCWhbVn72tgQvSqrasmhNhksaKSMjiwCMOhzI
pwFVsgrRg7XYaspImQS0TLL4kzUqaeOkdLKbqF4Fk39ebMyq/hzAkenVSB/vnZdCTNUqcrJVtCn7
6u3Qq+L23zo0jHnIy2A5ztuKVXLKnDiHDaMY7gNh6MfwOf93ab1fbR+NDDKoJKv66D5U4ZYN1sWq
/Q3ZvmjiEobfL6h78sjbacwbELgEu9qkqBaAAAQ4laOXS01CtI7tffyGCJIW5kMaVJLj0fpXrprO
c4Wk9hOWkh+/BgSWh/Xfmuu/0+IF5ZqvvFu8vDzwzdjF2h8+y8JlNeaphKX3QWVNEJge0f+fnyBO
N9TLIcta0zRaCTM04F2Zhhf9H+odDuVq1BRC6XBEYjjfTf0Apae/KxXaQAnAo950MMbnVea7lmKa
rTcnaTZ4j63w/fNHVYUlIxgwM+6dC7UBA5+vjiGhyMWJFcW74gJBbAii9q226khMrcEciTXk//7+
k7z5sdIROiPNPtEmTTxFaJ/Ud2McVqtceA9bYPUHfCq7xLbRi0E1rQLgFRg015LgVC4yfeqfyw+B
m6LmwxFoUqSBjIdLsp7KO+fu+s3HZ20vrQTyzoFYUR+IF9TIqp5gL0p281aPh2Gz9THQSQ6eKhOa
EyUczEcvYPOjfjuSfEbDmmqtF4AUH2C2kbMdYyGcOSfz/6MpPQAy9P4WrG03X8dpkIToyexsctoh
CTJ6GxAo1zZ0T7CaSN16TAoSwcXkPk5e3+NKIXboNVcS3wHQ0W+kFFUdYeE95NfhMt7PGhtcfoim
pBI6Pfg2IAc8jk/F3l2aMpAY1CUN1Wv2ChZwmleZc53A4sNNoj5tUGDkBbWhVaEATfTx37KdD0Zp
ETwdr3cAu/c/22MbWeJULodtdiPsY6/IZUJdwDQhRtX6lNwV/W4TJZ/OUAqAB3FGJasITSoY1mXX
xTPK7LqdoIP7OgVBePScr3AtIjGOKlvl2RyPPIpsIiiMO0ec6dYauvx7q1p0e7lvTr1P8ZwOa99q
uJ2/I1E6FpLMe6kFrGCsGgLxS1rWneGf6mZgSDN4XfnKx2AmoeRr1vwteKkGi9R68cXedSwEMJJB
v5ybbsc/MqcZMl9l+8jWaylzKQeXLZUJwdnEBHkGjaVqX3ahGAVt7a/6uxIeb5ilPTHrMsrG+LFl
xN8dEojpkK7prDcl/a2jZNRMiL75aOeEd//sOiUDYHqtJ2zcj8cCbWscxHJy+EUTF1JrnG5TVgQA
4g9a50utBaxAG9isXSHiPo8iE7aPoUvtotmb2ImBVm7Fcv57rwZdJ8JKdk9gq6o4l406OTGnNABe
sMMIujfQLNrCzDqfdhJISQlcQnoADtwNzo7YB+T+YCB/goE5DIJTVzgcPChROw3gj+GH8WHafZJH
8r7Hj3BOhN3gRxBZjXOmjIjDh+tktb+ik/aSwEu2x+m9p/uDa6RyNiZRjKOHy0E7vEgBiYwc5+uA
HJHAF7odMslx7IPpnIpcG/TeHWgUS989KWZNmBjQ0e66ifJO1bFhyMFvhvcj/YpC3O1UxlBzMxbx
8EdmcpnOXGT4abcaa7eeRyIPjgxzh0UpUYol+lgMENTsdu7dxpaUFw0BrIL7l9dYBUghNVIXCv3m
Z6AfJOYP3b6RQCy/LPxEF4FpPZJHxzgD1d254C7p8ko9Edj7FGShaOqm60KCRfRFO4QFrQU4CFMq
6VJ+XrxshkgtA2SDNQC4/2HfzPbu9VHQ8tSMtUHlSNKmMqwudPt5nijPD6n9dVPGNzW8ghXGRh9k
N1ex+/2ZEkh4gwDEjhIOl8Vg9JjRsKf/UMhPvOKyEIcaLIHuPzNx7Szo+SVVHtbr7ZKOix4kA1aK
iiICsIYRWtEmomjy4pfmJO4j5WKe5ocGR1zrD0GJFHwaL5WNZthYlKkrESHn2eZc1al7YLic5ksd
ShiQ3cwaPm3G/faTell4wEN8Cx73y3pGuo8eg7vN5hmPw+UOjTWEphJg9nhh6xLWHmK40VAAg3II
Eyt2bwjb9/N4guZuWD0lH3NSikCG1HcOKYdzjEm493ByCa++QSrhCHtUChfG9rSCldm33fdaWfN+
8FU888HdPwTHEWOpKrX/mRKO0yNXh6lJlhwjCsdG/ULkoEAE8mD3B3gLQ9pcMjCjDv/uBTCCDN5G
6ZswT69vDpjZX9/b76fbQ+dv0j36ZCX6TbpliQbhxnm5/Yq9+ulGVifX3dN2lnGaq0jmpg8KszMK
eZNyRUmzfrj19x7EuMjUi0h7ReanrDQsyQfeC0M3n3c2L3cyxoWEVrqhYXL7cqxEqpOMppXVjGPP
hmNoPT/lRRw6nlyPV0VRn45qfArNeMcF8gKEAIhUCjfgKF3oxufe1uTRkyYjYDbWkt/+/Xw4Fa9m
37Cx8+/YA38WOIgJ1PW3/PZhLryQo96vtEF6o/SMKf8OIe8ZNQD6hGy7QUEMCugASZ5nymzmGtKR
/oxy3huM3glWpRP/ShULqZn0AMXCp2uwQgaC7ai7pOVElog6jL0KoTP1Z/hlguIpzRTdZDuEnaQZ
OfJoerXL7P4nUT7at3phpeH8i7D5ghmv9k6f9ANsnDhi8Ll9Zu10opjPeJI6VOU15qm9hN7MrbaZ
RqbsDVA5COoHvkMc3riQup8VogxzdNAFRKIKfh9RgUxyMoPhmjjeurPHtX3CYMNzdNDz1AlVEjFk
IhsLQBLYAtPEFEwyxitKBFa0WJW2a6swhK9Uun1UVVfgxAuTU4BDfoqScU1xc0LCcBQecj4pwfap
ezQE2zU/toVDoX4qKTyycXECMfTi64BE30pROha6mUlVvOV/sY3MlJkP5KGpk1lJ37wNsQ35xCnt
OhEn3tmhl2zT1C7GeRGB1jbZllBL0teQyiXNT8J2N1uCpwhhgtRcSSKM41dbVO+n/YR/J4DbkFPY
1+b9B39oXXL5eKQTGRJIUTEjjt0UkIQ+TqgcPoVZ5hXSI4GP+Fh4IG5CQW1vunYhuSr3Wn4iJSyL
8vf5fROa5xcDLVHhtT0RhobigwoaPouhruwhpbUC+HaTf1hXOrsLGvcVjy+ThTSgv9eZjDXxMJV0
QdJumBPrd1KatP/q05ayUO6Y3n63AvLAheukETbKnIu7TlMPJM4vOz6WKMA6tGpOht+OB898mYot
+R9oSUy6RdbKRPu07kpPakdra7daEsvkV4kqRmBCAPQaw0HtUK2BfjDK7UELYWigPug6X0WHyrpR
cFjj68oyj6kJNflm0O0UGb8oc9WTftyROvrMSHGpa2MO01QTcVJHlfQgQWodeGBNwEnctuRMtiQ7
6AB04dwFdyEnUl65vbdco3WrWZJjGKu/HThgnGga8UEzm3ACBV+8BcBrfyPHtWQNMhco5Kw8EQKS
/J05B3aZR6gWJ9yfYC4bqUeEHXmseAqVsRB8FNyVtUZzZokpJT4uCxeOD/sWDoK0QJAJ1VlA5kVf
5HpRNSK5r6s+wfAjUiWr+nqjC6eSCkjQWVfRPc+RPht5FlqS3hk8S5t39hgR5At5B4kqYpU2c8ce
kOI8zbDOS93HbyHGmeWre4vQd9sHZ6RM7NgnpfoU3spvt0Pv2Uf+0HPRoYJJu/2tYbwiBBV+Wo9G
/csjmDkawut6gnSIjAJdFuuKG7IYQfLs00+YBZ63lormFjJ9bFSgYXLE1BB7476wEvpVVjVC703P
GjXc73pNQ8PYLIv2t2yUmSCHw0erKNHN9bUxQlNk4a16B5bhFN81yzlmHCPTiA0qbS+HjZ0lKkBw
P1GpvEgFKKTOwAyf5VcMOnXEGs/u3Fx7obdhHmFrCaaUkJ351lk2ueUJojtMkq984HGkpUhArcCu
yBP3fRmlrjSs/2MY09GyKgwRIIrhlbGkF1E9K0qIfyIg/af+IgqpWJhl5nip1lGIG+lM/alLHHeK
gc31+fXLwa6PTmC9eB/NQGGhjPxFM1sDL2SpWj9gX9hc5HGO3/uYBjlksLNUsOXGFAEg4ejiyU8R
rz5DEMoE8CHUhXftN9cFU3auWTzCox3diF+OAwgjIQ+lou+R2QYUjp4tra/yiTlVDBwN1slZDwLh
89coMMHyCndkKpTluYkvLPtDvDeW0SZm/HAuBZBORCW3bqqFXEWTOnlt9q1pBHuCQVlHjQtOsigD
4JTG4RWCBb0PtMa+DfGWdMecbvy6x1oxK0FVgsTnI1zreXOG2VoFMddqvZNAiGhdO3hv4N960/x+
JBJZhwEeJX0ZzUQDYeBjzo1cOdwddISJbR38ylCb1RdRZJg29kZ7t5lhXgTTbjBcUB0VbBkX2DUa
WyrT2nqpJqnArdo0qozDK89ottXM4eXi1HDEQx+WsVknFt2f3GFDRAJGYvaS4mblDRkG32wM+wnw
fxufWxQZKKa1EungXdqY+g9UargCVSqYP5GybNyFDA+VbQx/lkspWOnGtBMVmT9wNDUijvHbPqfg
hgLMwDhl7UFTzd4AnUnZqBislx9N6Ct+uQIFhRps3AhYvM5ol/x7iJSg98q/go/jbQT/HnH5y+9m
AVZ4vH4Ted4qA7CXTdASJdDDl2nh+6bA74NCQ97Luo+7UtH2e+ossTrP9s17k4oVhaU58KbpSk4A
LSyi6cf7P+puJNSF4uoAT/jwb8igvcHzjEimtQCnoefW4KyzbYKVHrDP979Q+Vc6KEaNeLNP9JBt
PfgQMDCXUx0iOq2BnCsvtfXHBzxx1lixTY9Ri4aOP6bnD3o3KegVLGfaLP7TywzqeoMFX17HXMVd
Yvzyc6uP9M86esj5kFDC3fDu/DtfH+mMC11HwD0FSOGcPt0kNfi8M/n3ahUbtjc4ytTKECeL85ln
LjAnVZNcovGruAioals/ckY2g/yDSRAvsQ4OfbQ4KLR2gxFdEeIiixqwvk2M2qmnGCQR4mCLPgee
tfKX61FAfmhpFIyW3G0s/cs0gurQaof6MbSLB4WamgnscTTh+/AB+3M0G48w9EUpEq7JycQl+cr2
oxeKciXa95Ot79NEFrBLeQXKghIIlz/sKAgtwVCBY51sng2JrZrthqY9NTDtiOpOXG+zOOASILPl
c0PiFXxcWHndZDt3wmT9io07jeRoucJwJ7asKaX5ieOe5zl+w0JN2e0EfphVnPk1B60n7QT+CR7D
xNCIwY2qWxHGWTE1vrNCzU8ErnHWnkLRDHXnn0X8GUc54M6mCQHp+fmLDmOVhOjQlDUynUIfqtpv
Ip/lqzajzW6SCeNZTbTZ9OTWvel1/XDx4dM+LQQDMBzngZE8X960si7yN3oDjf9J6/++//c3Xpjx
nVwet38nBTCrhH5e/bIsszErhX6xrnGIZpcdmozkToDH2NDk10eAfs68xiqCt3T+ku0RZFef2VSU
+YcwgTPM5l+i1nL6t+D/JUGW+M6D71erRj3t11riWL1wbFU4RDluNDllPuB0wg506Mz2bf6HhK15
skIoKbyeF1Sk5TnN+/Q1r+sUhfcsSjkj0jbYb3sBGGWvSv8SJYkzkHu95bGox8PlJl4MP42jEPnc
ok90nFc6FEe7vW3j2wVT78U9aZ8CI7bI1/GdRQCYGQ4UjT72pO2QNyL/s7AAYIHf/C5DixfpC6Cs
l+6aGCY16EUESQWSFc++ymA1Hw/2XTtqxM/l5FCxhc8KKef8L94Is57Y9ibYbP4rLtjyJDSf1SkI
prN458msd7PyCyci2OOi+itt0P1y0STHXsswChtKQP5nqt7VBVFBDXTTQ0CyWv+eQSjDjKL/S62Y
q7zFN0lHpeHSn1kgOmIgfa0aBV78xny/WmJse1ZwC0thw286ULl17NYoktSiP7893U11dlQza9QZ
7D71Y3p4jC4naUGgr6RVbdQS5kvMhZcCfHnG2UiAOLOnXEhgEuQNu7jfWgLSh9I2zjMgzpdBZiDj
RtgT/75qdXFhVzcNWGHYsNXWUTkg7/5+Ji698J+IkaaUcXCguYgqzu3JpajRgs4DMHOtQ/JA1uUM
Tper5FmKRHDza7xH9XfLyi2Dq3mE5oHzT01YvFfZzhfGXGHDFsbkCyuA88eSUY9wQoNub5wNTu1S
UpldmNjoNFEYEQLv4h2uVPUohfBdwc/3PnpSNmLDn6grVVurwv64BSlYf3olgVsr4i+M+wFK/p8M
eRUjGqcVXH4WMcOGdQkC/z43fnbbnwfmiD+bRmC194ALpmiQ8Kl7FcYpCYNtZpcWtxEdCwhUsliq
eBcbT8I6quy5+tftCg8uIfsf/5im9A5VRpmIrgPebX8o4S3fHTPTKqaCrj2dhPX7bSL6O8dde/Oc
iHBeYArdYhYMuws5UnrCYqFDd4rU/P6JnWBEKwO3yzw3NFaHxs1tlpPI7SCTl0kLcdKk1/Yo8XrT
hnN5tppy/s5Q9qiTlYgJXa2lVPDemjPLxGlR1Kxtd01fSp2Osi9pJuRvhQt9/V3CtuSK8b9sGiFq
qvBS1iKCVefSl2Prk1Iux3GfnNh93u8o3p/IcRoSDoo/7VOt5109aznu/1JXTl+I1TYz3+5nUmUd
yyouGzpJFhQaSFyVaztF7ad6X4l6gAout8TTCBm8JKwr+G5df98l6PrUMd44fV1kWcDsabLqfHru
BlzXFnoG0nX1KHP0u1vTtz8rdZ2+tYxn7fklgqafeiAg1iTHu3opq8BHKdDgRDXpxRjtj7tfqkpf
Xm9cmie8P6S6sx+921uTCfakgS5K8oik2bO2EJ5LvxXLDDBnh6UnGft35BVM/K69nsqnWaqw5nG3
78AAqYoLfHXiAFHI4kDZbN4HlRga9xeSyv4caWgkStuLt6H43HBtYdfjGj5eN3wX+XlT49zLDO9f
oHPXEtz0ZotFwOi1aOhDS+1aKmLubL6BBdZYDSEL3aHdnm9soEncvLKGF2qsYGwRcADBlZC0G9Ol
59ctv0G/engp7StVb5nuRtnF6kCDiwnq4ojwEeKyT3G74jRbhNhZ3pkbZGofywn28C2laMOPKyEL
T4R7XWVdnabyTkD/A17uflWEg6ZtUYwGDoOdAoWngRmmcPVB4/Tn6kkcvrZLaemYCNtYwRi82for
+TX/XzKeyVzAZdFSAck2D12YVVgSgB4GZ+PRM824yLXhfIK6ufXB8Z3q1HamqmKEfcMbXwN4vzTQ
+12ec6VNF0jayTS2bndD7pedDESfg0/V9wqYBQtQES8tDuxLD0akZFlD1MXduQAW+puqlWIJlFA8
N83WvB/aZ70CdfPTdoxtK88P7vH3611/flUjvFZZ3LamhViagalZNHeiseAZZk1NvEXsYAKReMdE
F4wydKzOZiF4HQxdvaHVLm9+ePjEzyyw62y5nOw9dVuxWxuROEAfIr36wiPdaye2bfzCMBP99Nhl
5cWM7oAShH0XkljMUs8Nsq8uqFqWoH56RTYMxlNRgO/lyke4JZ1IGYkuseZ5y4AGRrKjCehV3Enf
y3fXbXKKywwOT+jIBz0g5rHGAY9UXZm5Y5U+8aGDoKtIm3B9Y6X83kYf8uxnFI5A3OIBpMptKbyB
dQUrMxMsWxylr3QTNXmRcCuNHN42tXve2SzbIyeXvDczqQk1PTPtsr99WmLEvIaUnyDZwtWJw8RY
sBCjN5n/LYGpx83iqZ9SzlS65Z8qhm24nMAmOQYfwWaMQxJNTikm4/q79DdTRdihI8jqpw1yIKT+
a9JogmPiv8aqiUfPzPKy9t7vfqXdu12gWcd+59Pe4zJCx+02pRvPs9iXGbAf21uHgY6KFnma9hB2
/VhOhhMLMrBncEGRu6L9atZFREOqpox+n1nmnrxr5OoF23L7MkxvwUF2f2flzaVyV9zvaJV6sDoM
RP77HbnkREb/Dxw/bzty95pq2NQEfcyBFwC7FS9zPg45T8PqbcNdaMQoSHXJrwgmqlFWc0AlXJrt
tfDkuyUQJSOVaZJ7VKiZ1FVPc1kaUSswEQvstHqa7QijcsBsrLk7WXon7CmGEfNC5yBhZlttScDT
1y11zjesuHZb63xju6bDJpSvKiw2Qy2YBt8flJaJfhWqrsplT1tRLiw0VCqOn4wfgIhT7zGSkswC
wVwa7VmARrIDRAsPLViF7qvZXnC4DD2Ujs+br8ygXpst+qSI3C0uLvYy5o2yNSpEle2nLWEh1ifK
3L7j5QhI5hB8NhexMFUPSfdkUcV7mMhnN8mV/361PslXBdjDP24jEDO79ZLJhZ+wOvO4JE+bRq2z
f96ePaYVp7ovLt+3yjOiE+lutdAhHNC/cvxL/fWQof8UJMVlPDav4Mi1w/YSKVQMWkUq1J+nCDg/
glF80Yb1KAXdv7XH4mFOeDLv7q/KnGh5ceBZ/oTxB/ovY5jSj1WTWW6z5X7zgCaKyPryV7KWm3+B
CeAs/mWxm5ZkoTg/2bpqOoccZRJlFV8UYIqmxOK+uUwOc2PuLzQ4hkQVlt+2Pn/X8v1lf4jKs6BT
U3ERblAsFrkYipShut38XMJydxiilPBNI9hAXz9yk3Bkig9QXX1I/se7qGw0AhTnKaosJ3JEC76S
aMtUhJSOFewrJL7eiKT7nj8X+7Uo6Lw4yEhp69lu081n1k8efklf1MUyGt0OxFj2zgsfmycbZ5um
td92uzlF3ZUXHkDBrsai3e+bhUgULA7Imo/kNQqk5+tSTYD1z158zcqGwjuRLlZO0oeKX1bhZdZZ
xJDm3JA/C+RRETuVqBXsYZKdUp7Dm5VpOAu/0MTGJ2VL5oO8wcm9buRKXr0UBcL7HZ+kmwjxhU3G
aUoTPp2omAI1au0kcyE+I8QjidDQ3V5IoJXLQc2GaDSY4OPThvSCFdx3B3ERx8eSs0h6IVLPWCBa
9kdCYzBYCYjfCZ9tOorUb8Lapwo0gBD2fVtZG1snd6Mqsps+49zlNwiQAk5OOR1KQQD8U0I5GCbR
ubDJofWuuDjnzFkueIFczAd8z81vjV3Zk6lcP6txAJfK1JfEbbqZyCYNX0g5pbV89d7kLgiNZsPo
jnX4nlc+1F3t2LrT7IWy6VdcdgnBvGGndafFQM2fq58++0QU3n5w/Qxa74Kkqd0P1MYLIKQkqLq6
inwhDM44Hf/F/0yTP56EmSguWaI/lpwO4VG3oX/P/OnOgWBL2e+ETPenaI834Adf3V9QKYEa1uQ6
GEgTglBHCK59CArdPHliomCgD91/qcTN9fpodDvoIJjk6sVbZesEkr6mOrTW5RsI4nuMXLFFRUQq
uWF07m4VVealeRBHRKEsrhQzw2DiVvv5eVFnTEpICZjWZoTt1Bgnk3xQzmz9i/f83utwhTlw0v1q
89CFfwrF1DCsvqErSLJMcC20XF9MeVuT+mkhetpRxXAD3bkj8K5XgpNeVu7FbNWMOSNkiAXQPawL
iVOdwywpLrscgq5+jKiKE/6xFW+9egDCI02qNJaWzcWzzLWNznbzHXVt93m7qdwCCPt5kALC1BG9
fjut3zwg+y3RhYzX5S2QV+fy/orLMmh++P0AURZZqguoHJafM/bIwXw29i2AWIQy9M84X2/A3frz
FDh4/30+AULJPYnh2GgnIXwL7t6LG0jdfA+WFiMKlGDCuf+u+zKHj1olAIM7Iyi9yDSgTJhQd/OF
ZP6LMPZR/8AwDHnY22Vsw4T+NmS23Ene8DCQUTMm3169ZGUFS50NmfZ+n+Rw4Gfj+FYFql1me8tE
ZKzB9OXcz4QWRrDeGdI1r8KnofDU/jpfnmC3aBAoKDDz6gv2qp5e3WB9Ui+0gmNkpzlU9XuU73sb
Ct+oXf9gTQKidJrFxJv9x5eUqk5NLWMHcgMWT2sOX0gfN1WX0CM5uBEJtwoXWkudtTkfAGumCN57
CeKwYvCJls1jnU3as4aFaPcbsa1jrjkS9yGzBOhHbXD9XBeqIUsjtH6SZUn3NXNmfjdLsD2jRfBl
4usnud/Uhngisd46ciVzxb4BnP94msOzZO7JpbFCG/Yd6exEZup8+xTfw1vkr4Xhdg+24TpDthfX
NnA2U13QOAW60prGxT2qzNeYzpf13Mclu+oRcRUs/r5NWE1AKyYdNeg5/E5zciijJQiyZTTESAn/
WhF9DVCsS2pgsDXEf+z8xWMnAiB386fnv9W4AlpcN+pM7/glDqg6AcmUjSvzsLaGXTovjTHod68q
8kmFitk656p7ZB7oxfQIT8NIcHs1sBjllC4qV7S6nX1ojv+w9FS9LWbJdiQ70Bczz+oz51ZstqFx
xuT3USlHDsKZJVJvC9AlEz4s6vcpFLNc16KbF6mHQr9TQhe+L+hrW2/1NXwA9fr52ZtXyG4snV1U
+pPC9DyKYcg+D2zXeuvzZ/UAjsgutPUr6PMas2IcyMPoWsYhkU+5t0XtqVk4xrDOazr8XSwM4sfq
JGbjuI1NznOeWR4lu88UCtV04rHIh6csawM2bDzuPCRt52297xZO/n3JRtLiF8Q+e6e8ksVN6cQz
dTOlKFLBGVa/Q2qgBQEPzBi59ot5pPyhN0izVxUcr+af1yuAYfK/XUArZe1Mv1HJRToXq5K5vreI
GcBCn3ZQL8hNHNK3UUl6mCFy+YqbDakSjWHYUlx7HYramRd7YpvD+SftEWfFD2V9pcZe/+Mwa4Cx
Jtlux3qk9pszhut7Wh2AN+TZIVikkGfjfVFGVRneZda8jZIp8nxJMPtVOueaqT6s3rTFjr3wPFLP
P4PTPdd68wSRXCBd2t/IMO6z1PoMVs9F4dmlZW5V6fpMhbL2Y/2zjgMYoqECidhgJOiQ2f6fmv4U
m5L4JZpSNzGf4UVb2PFrwmnamREIrM8BOSYgYbzmqRZlwpSC+qrIEEcaPz67W+hkxCewONeKLpV6
IEvSphDG0WmZYshbluA5xVPaOpGw26BsOjvYMPjsijhFaPhkLci9feFVzsWgW/i+I5umqlTCdMrz
ErRTRFhT5Xvnh49tW+x7WkqP4ihAkkrVnW8rACyoGRl6FylHrvbKGlIYa6cHEIvqLeoyyKbLGjnB
ls4QHLl+EIJ7+DKA3NIRLFlH5UCvM5GGDfekFRD1nQlQTbf7qxLyeadMG1e4opcMHkvOsHsJ4Qnx
hkWlEvW9j1wqixjJseqPp6tJqfgfsyuDa7dftvs/ENs/hgfbe9iXyrr/fmNBu8y3+1t/5JvWuLIa
355550YwHr7eckVzwGAdKO2EWP1GZzzh0HD8wbK+uhAM8TlwF0zc4Wm1fviFe6C36ujEUu0gBVIS
fdfZFVhrERy2rhw+UcEIDxdBMUjT/ZTXLGVyV9JKtP5xfdrACDEZqDUczsoD6EnVx6mYQnLI4wzN
DsZy8cWl8+wGfMA0+XPeO9aDHy7g//ED/jq+prZP610VhtaYQD6abeXBpC5gNK8iuITCw2V+XGNc
Wtx9ZpJw/WOwobXZQ0mzD5JiU5bySuxvly52GykSsnmx3fBDw3Fbxz9VGyfTJD3DjQv8haJDFgDw
abQeIYeZMHxQCXoHMLJfvZx0iXW22kz8FzOpBGc5qpIqCAD5d/0W44KJn7g/XN5A+/ZuzmOjqXB8
fTXxamV0o8+QzQ1K6+X93qlbBx8Rd3X5XmKiZ2RrvUH3R/iFzg3ciAD9IoVMSSzAuw3G/vgl4g61
t2hYswVH1p7LJxORGGn4iCRnvPjd70bg+/DTaQo+AI2XxDpb3752wej06V47jUAuUFbQBv8fmZl8
d1WojkEmf9pwmQ6Y8Vit93CfEgQPFXBgS7cihu3mLP32XWlCdCBtMnC2Uv1TbZy+fIOvQ8uNDyzj
8MTc9eUSrHUAeqd0mQUWgsovG3fTevZZXe9iZpjc9mtt5UN0ShzbeU89J4GfIfi9skrQc4hMRlol
+Er9DZiy9AktGixdzUZjnWuQFWezcVhfNH/+dklaXZiQ1DiPUfxSda4imXD836pzuF0T88oOiCC1
+HnAEJkY/yUr7qE4Qd2/mW5RKzaafwvF++AD0lgOf2I2sTjn6XrSyxm1gwaa87hps1ZO3ZiJHcaH
bGLsaW8aUTmzf9FsaZ30/niIzEuuGL4Zs5Pf9pQfLsjRrQ9KTDqEwhiP30iaxfw5Efx/YuNP/L8v
TUW3VzCagx9yXZYL6rirTqwAnM6e/QUY7krxUDgPoG8IDfKMY3uHhyCniP50mQ4tfdZjtZ8BJMNm
V5NEPXwwyoeh9qnJBMGGkAwc11O4YJee3v4KPlX40/7BKe8bWG6DgFz+f0JBsiupTLxUnLPg4/3X
UFaonAMGIP24v846s5t6/0QAskcgNzfdMzJtwuZjF7gsbwLAe3M1wY6xtAsAu+a//UuTQJiPS5Yn
l/SU0KlmfH2/C7B8pMk6b4RC1L23lbpjOOiXaHGg97qDtuEPD3ULZvWSsXij9ZJ3np7/X5zLxox+
XX/U71/K8vVQ/WpXfms2OcXY6OuHxI2YrMJGoTX+6JSXjJh0wpBucvH3NRch1MZtrrOg2wO/juII
J02ikq37qcFWoS2WFxyMCrEZk5iPUeWPMn0XhvSV8nKqYCzVtrDbWhGa/8gWIqwLAcacMUNUVQga
TBSOAdPb/mEU6edHZnD/qvsHKEnxFlh8JZmC54i+bpO3kJXpwvnFBeER+pS3ND/5K97OD/WiHgOl
E64k0RTXaHwgNR4xdW1444VmoHFo9mJQa9Ewh9PKZ+l8xt8eqHwS55xm2xDJ4itBB3sfJ/3V8T27
zanoRJf/UQB9mu+LTY9TiWhGQMerTein/tgMUDaba+cLhVFqy4PYfpjuhjDi6tJXgQmXl3Tz3Uvs
vVeADLE5/D4SdLV0V3xoQf2fhnphlvD+LTwJu828Y7XAjLw5a4AFzxXC69pc/cwG0S/J9C6jeAKv
aaD5o60qUeuYYYRvZWGLBlAnwSopHG2JBhaBxdInumY9JmQo9BDGg86ekaBiORMidSw/cahzyVqv
Z73kDp8F0yusVa3NywZqF90g/YNxod738JteD88UDrxjdR0X33KV27WmdhfU1XXVIIXpaulAd2be
3pqp+rPbdWo6AftbP+KishzTzCqCleraWsyaqW7+PIH/qik6SfQjQRCU6VpOfxhcSmYSYC5XZmUQ
hgIAiwy50STcZAgTwqnnkjb2XWrGhAzjib1e76T4D3DEATwm4u+BAsYZsGEcv4mEe6shyVrl/dTg
RgYU7W1mxd1jAxPJ96Fn6y2GZHx3NWE6d2vwYw3pNOF+z9UpHZde8SQpHVIkyfy/beU1LJLRHuYl
DEB7YkAraZGUhZquyUoyFdaSGXAatmVaPrsFVJbnkN3pXJL0qsBozSFJGy1RE9TTYA0WqbPRoxJi
y8Z2rDpvfz1C42g/DME+kPwXaz1j4bpD7OLs0/Ru7TK9lop/zu2H3gM9Hy202sZMdAIgLO1NhGXB
XatwdMiNY+lUw9ohguUvOkRnX0Ae5tTyPdTwiiwEm6kAF8N1CRvcj/KyGM//pQcLXTHpczRu5i9t
OJw87DsN9sYV6WgVDW0pHvvRhp2ArByy5QHnJ79fgWA8hmjM9snCN21ntpPBaZx6goc/y3O0bZPX
bJ04f56EHo6quQNk536xoM0F9ex+vM0X6IFxHwr/4D1rn51sN4XZWn4OQfgjroS+C6TRuzQRkIca
eqB+81a1bSot6r0wGjmnxtAEPMwMdGfec68RzGjWwK3o8sdXpwdfE5zo5tzXzjKgPBCi1KAv78vN
ifpEPxMCT1gviBatvTHT+kGLymdFE7OQuWEcXP/kp1AIcQa7LVJrjL3BugrY/eJbVdL5nHnohAh2
6EG+HJwd5hP6GMa3m4frbITZ2tokIH8LVOsvlPPmkGa9PkPHORVB7WjKfrMAyVb6yEhhstfwpmdH
xbXiNibeaA5hjI0IevV/ak82xd/e2FOCfIObUp02cEt/0V358oVRewlqy8h0sTaPxTEawk9z0lWl
JxjTf5pxuj6y/KBuXG7fO67se2LeC1XIXNS6XO11HZGyjKqUEcMLp+Sbh/o/kuE9z8bND/Lr69N9
rh87HwuxaKBv+yPm2sDBLvn1+5branrqm931BF08bW/OGuBPJJw1JxLM6B+ggjs0iDbXnwQqfWk7
//REhqPr7GwGAYBR3GTSOASbUIVndRBnOPKt/g/cU8a+DRdX3Kn4VQ0zNf8QV0cgUKJCvNrJZCXD
uRR+zsLAhe+a5LM03+hHsoItrUT8TDunxcRZ0nc+Z4q+lkEo2taVbkBpGm/QV6swIpZ++hU4KG0o
cYDP+eDlG1aJst+8to1NzG2M66WlNRCtahkLNBPlizQAAnEaouLFMqHUlOu/yrN8xVMg7jZOh9fC
+/lUnD/Gd8bflPnKRvPeH3ziH2IlYtQvigY+OAo1bS64+QRsUf77NAR8I0pxScTF7ozDgYhgcP2C
pYWy8KWMQ3qN+gKX5o4iTIzZz7SFwSp58ZVcvN+EsbHht3VH405r39lDWbTIx695ea33oshzw8K7
jDYvoYCGMgM7plxri/rABhImvPKX3PhCwbKRxPFOnblPUa7kSIi6T3O51K62VA+LYEkSB1U8e+2e
nLw0nvunTDYUpCeS8gOdAqCtAttUEn56gcxUVeN//XHUq5WPauogLXMMCmvdWoZo1xv2ifZboO9d
IBW8jdI8FkuUX+MLWpktofQnxl2eYmXT9VzYt3tY95gXWy+8vNa2scD6wnUXxcnmORWIGYcRGYkE
DrATkCXxKSV4u0mg29CR1U7aCxUfgkY6S6bPn49Rif+ETDJLDXOAMczN1T8iQnFbtidoJVe3Jp5u
ll/OApeegs0kjkqaGPMgDnbMjLcQxdb1k5JnrUVAXlhaHJjbeYkjNND5Gq4/1mYVgCYe+wTvuikh
Z9Zi15q56O3A7UazGhfoz8hQcWkhmEEhNNW8+VHpg98GLSK6FkPUj9R4PRxWk1ajQmfePodXAqPz
QUSlvFczVtP/709UkaKimpb/i58uwvnkUNDJMezwyONinCm8klYc/Db/7/UWCOOGN9pfiUZh09g2
EUslckDvCIgBFvvURqOX8/ZqyiQ/OuEuSdUIpRPb90dFTdbGBeiddLA1xuQcFcrRV+a5qNyApwj+
f26mfLG8ASYRYvex3gWcYa+qIq99G8Y+zvem8122OVxZ6bfAfftZliYdQvrdZhpacy/97m4LZXkl
eyj2WwKcgoKQN5kycU7/o4n3U4XflU/4lNWMn0bgNzsKu+omVAGscF5ViIdmK11gnUAPGAnRQCJC
bu7Fkm98Mk4ndMKKc6t33WwdzP+X/m3sNBt00yRX1uNOomBP2HXpkD5WC6+CvHGcIxwMZWYS2h/W
pHZxb1inOGALEdeVj0lSA1zyNN7Y8/krGuvDp4fc3FXEuHHsNbg+aoobzBiABNm26ZBjhwmzEzfU
dqEGnMkm+oqxSGVMh6B8q7kAvp3+xLgowPlM877MWE0WXulQeH757/dQy/XIpuJo/3ruZ6VE1zMN
GKnctGWwnIwAtG7AoYcUSfP4U44IncMeWD4ljNdzFiGYrGZIAPRm66v40IaKnWOpllM9FEQrdLf3
x0uKxE4QmT6+WxA4nBF0TOvv+B6dhFhjYlGiuMx6h71mzcy3nYWb6TLEk7agvkUAXuUnNin3vFdy
PWPvY9q+Znqc6Irnp1OyILo+Tcgo6MePn4XEGLDf30PfnwdEtXf76752R8v+toQcWzZC+dBwH15v
vuzr5W4rZ9ogxbOs6lhjTuuuTFZ8p6Vsc5JkFsKF5l6Trt/uqAOcUCoCO5fyJFNVN2JQWQtmBtiy
tLzcUPeG5Q733f24DDHbU2yKI5jm8rvBtYtSRAg8xZjI+s48R/t+9qCD7zWwLzfQPo7lpAzt3Ozm
LFzUaMkpl6UsV2RuyuYxm3C5/zB1ERQRGI6NYZQA9+y5tADjezC57XOBVqFlecxUa3u7OMBG1ds1
CIRX/wvg9nQuCux0+4FxDhm/V7mCzL5h8KgM3FUD3cKPFs3ISHJVXDpD65Amv9Z3mUgVhNB/VEyH
vU0W1zjdEMVl9K7OQZDPGDCN1h8kGSW8xbFTlnVHrQ==

`pragma protect end_protected
endmodule
