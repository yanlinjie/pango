//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2014 PANGO MICROSYSTEMS, INC
// ALL RIGHTS REVERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//the compare_256b module, which is compare the 256 bits data 

module ips_dbc_compare_256b_v1_0(
input clk,
input rstn,
input [255:0] dina,
input [255:0] dinb,
output reg result_equal_to,
output reg result_larger_than
); //3 clock cycles latency

`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="default"
`pragma protect author_info="default"
`pragma protect encrypt_agent="Synplify encryptP1735.pl"
`pragma protect encrypt_agent_info="Synplify encryptP1735.pl Version 1.1"

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Synplicity", key_keyname="SYNP15_1", key_method="rsa"
`pragma protect key_block
IZnukXin8r99hGPbiX7vaCNWCNnFnAld4m+9JAodN534IHVB6E5ZAX1BvcmnrsfOAhof426pEPPK
VM/ck+OsIinWRtZQf9wn+WiFtz2kZLbBIfl/6CBbEpOOjD3WkYFT9ubkDKlZkNV4RHDh5n7Ln5aT
Uud5pW5kRlAZ9Ns1hwos5ycay5NjBEenRwjZLbAb+k+ZmMYq8lWUMxQIoLYaxgkxWCSS5WwnB9NS
rXlUaaaMso7FK6I/ynEN40xSCMrX7qF8aNdxSXYuQ3VbicwhQbHJSMW15M8fqyIwDyQzvYvsk9Vm
GBz4Q5R3Uqs+f8jxt9mttb/OFQvT2KuVT6bTMw==

`pragma protect encoding=(enctype="base64", line_length=76, bytes=256)
`pragma protect key_keyowner="Pango Microsystems", key_keyname="PANGO_V1.1", key_method="rsa"
`pragma protect key_block
fpejrTsJ3J8tlKwtYHrxaUnIVhqu5wODIuQLgOq6eT6eV53KYZHTKZeIXy2CZaRn2XfCN7DZblA8
HgqTMJBGdXrrHKx4F2evDi4G04yWDjvkdt6IrvxRRzrRWT8XovbR5/+H9gKn0q+bK3yq2vDU4V86
gK5bj9cTslhZXHfUn0jv+0M87lgCColUjjCLhZOAqMULIj5ABirXfzPO1IshH7nBVlF7PGqPShfB
XDEcYW6Aejbmq8TK4byZaJrE94QB5E2coZPIDB7wDrh9COCQSoBjgK4IGvJSXkvHB08NDaMM4/Bn
qje52t9vuvAHiKD0Vr3pcbG7DcXjcjA1OYoMvQ==

`pragma protect data_method="aes128-cbc"
`pragma protect encoding=(enctype="base64", line_length=76, bytes=14000)
`pragma protect data_block
Q8O87MVwMoPkBq3TFn3ibJRZIOr8Zur6jxKj+UGoewBhAGmTjczMLRar2KZX4bPB+CPcEnpYoGga
oaSuDLSs1ZNU04wHABp+6j+uwIlbARgP27ak18heAQC9dmG5RSCwI6pkqWdlmVDu32ECKyv6fqQj
9MBI+X+zkcDXDgXt6CZfZYDnMF0UyQd7Fk2NlaUYf9O9CClZmU0pkKKdHVQchB3Q/IuzPHjSusPH
2yciS+eZ72sZmiG+m7fc24qFpXzIzd7G4NQkX7AwvT19H6eDj2sdMcPZ3k2EDbFrobro+xmVZF92
jmMBXsG+d4WGZauxWE3Wj6EJP1UHxazbAeZiY2jpef685IpO4aDHBmp68y10JDaVJIbft6E8a1QE
4+HrlbMdKq7xoJW++W8VFM/X8+9ej0iwgSgKOwsQr/JseqlQOXjlM9ZSJ2hVEaUVkTXhVg0YHqQc
7RfKUsEBfxfqVqHxGpBui+QJoJLexP7hKg3Y9zY/AQrbe0Fx83t+1Q7a+qEgy0+ozIz2GIgsK9Zm
p8aFajE03aPOxyZFOs9wS02LzgKzpOFOGU2LCuchymmAuY4all/7cC+COjDRmnMnzpbA/DnATGgh
EaI2zPuycQFMmABwENvQOvFy6OtVXPwnadTgYG5F5yQL+++oq0kF2ueuvNXWXytOU1/fL8y9lfep
Y5gO7isKb7lgO9Xw513rRwZn4v9q7N0Hf2jJmVy3e2gwE1gxzP4/DAQ9UyG3ZcJ8BZk24BGm1KdN
5w7yM0wmbR4ttmKw9n7LbrioesvE50J9vdfmEYyI8koOnklxKmOX3QqsX84jgTzc/7cNZQ58THFw
b6NqrtoxCwaRXIbRwX6/zQqrC3Zs5Qwlup2owobvto4Y6toJ0QgCk+pnNA9JiD9pdo3pEWiQL6Rr
CvSs8TGr3thoEfaG7Oe/5oYFn0yOBjb+O3dqGdKoT7gdkuzZo3F6le26r1X75+qL3fBbS0MnEmQF
c9SlxR6fNDKt2aIQSU6JdmnBT3exv0cHGoCFNnFyz8Oa7aRN6pM1g21zy1TnKt7muYcUR99zxVRs
/BPAX0W8HI6GR86Dy1oPuftMrxsKpjNiFScHc/3XapEs8uoTMWSILZJbFy+E29MXmYmgtUUgSmPU
YFuHiYgK5HAyIFi/nYOrpyrivo26yxB5MI05L+ChipU2FZxSyA3GmlA884pUeSDvVRxwej/ntelC
RGCrl7Kc3390o5tDqVMXeQw2rOZ1urBQL0uEmICplrmFQ46AHjmBCSAUfPg0oKA08DyoTFXBlebK
s7z/sFAsRMRv28BstnyZo6E74whv94nnk8SNOpodGCBwimTY3hZE+EunzO9nwIIhLAloOFP97k3e
daV5VTdeNBiKq4STVHfaQwR08ZgBbrfiLWj1HQw5NaArIQhxy46RNlbpCnCr1nrVCJIpzE6Oqc6F
bACDA7LYspQ32s2lsdoD/oQ4ixiIy1RpogRD6HNDKQCM/oB0pgSVkmXT8Mi0LZTDTA3hJTBe0TSD
M9yQSxP73O8PUH1bYjHB+eDk9XIVYFU9WpiRryIYjWeUNc06q+YljqYERhx/P3QeX1mKswiB98Yu
X59tsygUEbYX9xyNSPgRunEdyHJqVYBAou3Pl3WNn5HU7B6TEwwlMnK9JwD1CY6HxF21zjFIW+mC
/umVv24/DFc3OFF8dONG6042d8uCYBDKcMKReOFZNCJ3pC0lklJ50H44Xl4Hf6tYKJzt0CvEMwEF
2dW5ZfphSUuM+O8tEcVfNpLgAmHDRnNtWZY5ruhfvigRAf4WtEFwWBdA1pIRR3pSe9iOljiwvxGd
YTHg8gtNTUcI1uuZAEJCJB25AWd9KnA6bOFceRQpyLXrtskM1/JLg2z35+KlWUjAJJJwVERiNo0B
ih7PhlYs6Z9/KB9ewjYmpXOer8exqq9VA0B1lwWjfuz4UEQoVl4Wnr0gH0CuL6y0HouKp1h2UCNt
MNZ7nu9X8l+6qK8Ttl6JJhXoMG2fkHTycLhNnRQy4AG2fps7nxjQieOzc12QxbGY6hnNhQAGLNA/
T/uqDmIv7/1TN/qnK1vFerZNKUlsXYDgSAAsOoz02OHQ3/yZcd59RGAyL7BgJmv/BCFBZW1swgYM
/Xfgblz9pbDMmL0nOulrz+H9HIp/HNn8i5nYGogDRi3AhNSl02Op9BfUTTa6OqEzw1rN/r23dPTt
6ajHXWyvO9V/4eLUkHBcVXijKolFo3i3wWejYm1IlpSBr3Mu7yAELFERe+OsqJGq7mwDLFK6dIx4
o74q6GQGwjtIpUwRmBav6agicFu7dlKs04t0cAXF2wVPgJ2YSnaMdnfKutT2KsPvQ5n5jl4qvOSL
RAHbvNtCjsjvlVW8bq/KfYLvFVnoGeBMeJnOtOUHMrwnOoUg8l2wD/pSQE2J3btmZ83aG1dF4YP7
jo9g02L2Sq1LpOmWjdfFWPDxtyh6e0EhU24rb3RClctPtWkAoztVC8O7AWlD1FOjOkdemcTslByI
HhDWthupdq0pmZ+BKm7Q36+HoexrDwQnikMmpLuiZFAPhTTK/J2qnkZvyRgmgmuJ8sxqz5XwYnww
zebuqGAs94mJoEePeswjagU9MjVnGQYcpizM/KlNsnqgJ8i8LpgCBSo8PtHD2bIOE8+Ru/yzX4MK
Hx33pSZu0sWDHe4dqcjL9ljj/peixk9Py0jdpfF45K/gi2DWGUwGAhIxomOdMidf4Ro2d2oQPjLl
+Qa+TsO5PvWHO6nVKyER6L/C7zpFmAbkAkAQ3+iF/b+KVJxn3xT9HBwfSxdqFgy4ph8JkOwG8o5H
T6Wvm5xSLDACuOrJD1ggfzrlakvsVffnyWly0rkPIwNYj/lvA3iRds88Ryg86aQkbY8JIOthPotE
UQYprA6zktdxKrlk7om3zrXWktGwqX+FLSEV1vXGIEcUQNdDeJLi5wurhJP52pbEn2a1PnB9M8pF
TJTc+PQ+7CjeVD5rNgFgUzFlFCmhs5LBYlxzy6LQw4xKnKS/SSXicOsGGbUqDG6PTwwU/ZePZQN/
4oxc/yzl99SYZ1WrFSK0fgYI2/I2q8pucXyMlQdTge5tyF5Ue4ArARAVrtDnh1WyVupj79A9g+DT
O5fB0cyLDIdavxKlP5u00lq3otRmNWbqzqASGOtr6lbf2hw69dLrO6zT78D9E3lvJn2og8mv3Nda
GORDjLI5erZRpbXEFOKiiIq2krMBnHzwdD0ykJ6Xa0ZjHnXfuKqNwivEB74nYzHg5vHzi4TaZsyN
oWQaNSRCyZxlng739PqBdekR0Nzzm2tLHt/21CEnHePjKwoCCJhOKZd8/9x3flH4CanZPClpH2wo
7oU3g/ozNJVsKWJKOvQWhDCxLQE77tOzFKzzWIUCk85rmtsmn6ESS+OtGUapnFuOoaeLef5dwnYD
F76qei0M33QIIrWuC9Eo64qCRL4SxB6fWkYVzClO8AwM65P6xOGC8lehDdwnggYePlTGCGDGODo6
zAe499pxOohxfDWJNNmZ4h9ZV2bHboCSzpmmK933Bl4vo7LTC8x8J/ZXI1PXkfY6fEfcok9KRr2h
tnr8WPCIQdddW+Ml9ZfxbYNqqQc49EpMiEN5S+SScsjpWMbr8cSQtWNk6LcB6t078xieJnnxqLEK
sYnDmbUTneaXhkje93VQKXoYmR5XergppnuIXx9VgQw8rnxK907xsy7WzQF54YrR3KQRIBiugmWB
gcsTzOsrJ51HD70FLNKlVaRiypZfKZOuisOzh2StDcPjKuf8yzxSTkOvBGypM97ZcmF+SHmkZbGN
PcpcYDX5D52asA5akGTbTXMKB1po8PPjnnFKiZKOgga9AwbWXRScZkPSZ+iBRda4qBmJ5iQxlkte
gOq2pysU8mHVsXXfWOkmcyXpWB4UY5aWOXrvSDHyxNmMbvwRD1L1hhms860kUa/F73i6oBwtZHzF
EYS6otwbJm18IyKyv30Ock4T5MVqslG+8lwrs7vLQL34CSJl+GPd3/g81kG3D+v3rKoBeOVmSC3o
qy9dVAgp9rmipMvGoAUpVeZn6g9wGail2ip1aLtUQmSPpy6tkIPaX9JpvUQvHpRwTKehIFOg6JqE
kugQejKLv+E9pt7IRw7v99voob7OBj+9If9PImxp+ZODF15avGE4RiDhhFz8Q3tjp7wKRHxCqQnX
rN92eDsVlihp/FKQRT9i9gDZlUlktTF3KL23Pbx4P0+Xl0iSQIbz+WDwmb6aMi4t0znEmacrY1Kv
uCXN+0akFCVLofhtjfax1bTvneD6cnOcZ9h0mTybMgAwAiewyvCyzg3PXH8OZztQcKaKdp5HAh5V
0yRzlBBD60g1fAp9jo6luuLPhAxVfdq8cO7viHn2FDkOghtvHDnhy5qd+6nVm5AS5f6NBSzeRM4f
JfbsKo16eLqDWtdt7DH11fTHlnjmjUHJhIqUax+ZPNL146Bdo+LDMLZ50Je9GYjPb7oKiiovtUTB
CjYQYsvgnSacDin7FHlgxMvQiMpRNPvxoRwI8kEvkcghLiFcX+DhFlihQm1Kh148ZwZSm9mrPK3j
hyVraTVxI70Ddd76S3ZLPw+8e2mQAleLHkREvhNokTrvByB1jxHGkfF0/xSjNNYcNAMb7B5HwjMu
AcBswXCL2Nmlea0jD4vMAKPF5M4WP0FksGkphB7Zpjj9jVugCxX652qK1Xj7dcwPAp0rJfdmmyzR
BJayFelN+UXWBQlF3+ZgR1pvA1/DmUuz5AvVWRsBcPjsLF/J/MUEhDFzPC0HgicaOkqQK/SbH0xi
zlyvEXpqkB4EFk/zMTNjt9zIXyrU3Go4C8MM5vdJ27ZFBjzEWsuMgK0CNB3vYOTZcgMW63zZHTru
vN3mza0UoUi4PKpSlCWmhuINFH0eVh6BUS+0szwmE6utM/3/faN4HWfvbqLIurRAVxjTddN+Iw8m
mE6cWhHEhhzkKBMQCTrPU84Su1NGMo/J43x+dMztCsYjSJNORkVE/0s73jrjRZ55y9Tsjgs6g6iS
6wQalQFsrLVrCsVDPXH+hcf0ONUcOq2G08MuCyV2TpqyGYY/q6UG9aJ7jDyLbnM7epY07Vnu0DW1
/pkH7UfNCQmLUFA+NOGKHJxGX90Tw0/tycXm0WvZYgKH77y5T3DkquiTt70j++FeLB13LGUwfiBc
cOjm5vM9W+fJwN57wBtpPbPhC/5RdN7CjOkcHhnN25EU8DxwVwRV4+MwmmkU4dqUZgGKKmdQb2wT
ZMLXqDuYYw61blDVgFRElRmiffbiQ7eB5onuArgiQMsj5yK/fHtGhx3N8IICRi+dy+Gq+pnobAQv
YYQm/tpAcj2q6v02tKhfKCHpNbkxRq1rEGe3JA3M5nRoQmg2Lb1MiTTrG3RrHxupuo/rU93YB8iK
HGsh5cwbqznjnz7mEEdDFzbHK+pcbj003s0h6k4634og4vfBDFCZXKpqfXrleDQOHTcbcqBVaceq
zh+eSV7n7yjkmDw8WkXh3FBB1oLph6XnZyYv7VoSWIJF1XKa+dxBmsmP5Alvp+JbqgER81qw0kuv
lKxnv6e2ZSwBzDN7MAjN+Sz3C2cdi7S7yKj/HaGexpyPOD0yKCjMq1zN6ji+M5GIrFWEpM+K09l7
Npdu71JMBlXdn1ltQZ29/LnXwXCK3/Q5eli1gL6pLwXB6EYC4Fi2GqcxyHcEkZ2wApiyzldHnyij
Tku7jAptTes42gbnDbADPcyfy77Nl0HewBIlB8BhVdyyaQY/h1wswfCtAKCd3SGCa5QspkYY9Eg6
jqMY/9i+viMGp1DsMPjegc9K1JX/DSREM6tLU+vUgBlAAukmBqDuDjbTUJY8WNTqm9C73ni1Zb1j
z9iWqqid+Xh7pNwe2oKD0ZknXT8KouEkGndqc9O+SnKR9FCqyM1Wg9L3+g6R/M/ZYGIkaBgMF5Rg
T+kpkR/Lp1BTsFOzIYemyGF00AciGe9UnytayMzj/8miA90O/pvxsUrAaWukDtC7ykl9dR6xk3EY
O53J0DvG/iEJ0vW+X3KYb4DXt9RUyW7wD4EHXaq16+XweH9VqMTMXutksX2oU0ay+oY+FnFU0T2P
lokDXqKzeb9dS8yyatNDVNHK1S8rhrFjn2oN+KA3FRJaTn2YnSvHesSw85bti+3Z1Us5fi9E3gON
Y0HJELvmzxcKvFjgKnSsog3M3JSC5BU9PFjBrluKn8CHAUF6eGOS74MgeeFj1cBQkY9JB/JkLdyn
ql8UBSsmdI07Pi0efwqCF6+0HvgYchbzFFASFobbOxniVGPyOP+X2TbCr+ufJ2eHlNd8v8gt3qce
TBO3ipr7dyUzaDEBwANvRzWNkQt5g/q5W1t5gNd96Qte/iH3JNdOqxr292nlIixWLBs2GQjzAhEa
eBLTttXmUWT54U9PUI0rZUNVJUzHcAq8+EDBZmyecbGwPApcnVoJ2Oo3LuLjj26L/ecybZMlB78+
IK9OAykCWx+aJAfJfmkB01Bq6x7HPCY3NtZv30qxEuV/PFPyCez8dDrH4VhkvTlvgh1ew8Nc6m4X
42zeTPbIUqSzHvdEE3G5HpDcRw980M9v8zUi9AhxHSs7yWyTSdm1JbLwNJCbZZiJr10fYn5xofQ6
+YgmgD7XaPjIeddMf3RqH0sKqAOvTRWI8D1tK2p7UXYijn+lA/nObx7ohV9U6UKTG/MPEStIVP4z
mhct6Qw1C5Qd2TBsHshe8H3s3MctfI3SIuG/FPMw54KIDhQgE4zTBZReHFmjVxfAN0wPDyX7bHaM
JKJiGooxnL0g23xk8nD9P4zW5ljycsjDw6I1r3adXkgy+d+eIShh18G6LdWY23J2JezJUxm0UQ7e
WpTiMAXo0ypueqi3ApXAK5WXLTzmKoFDr7W4rPbq6NobGnSKMFpoYXuAm7gjCP0SWTTnng89WDGA
0YXUrjJVu6UOvULV5fS1h86JXteH3MQhgo4007JZGnvFh6xB/kpiPG59hv3AnpCkn9RxpNaBz+5G
ae8qoLQfBSXfsAc2rDpYCANnLPPTbH6DwkdwHTt5evgAYdXcUcyv4uDgNtNt2s9+ZuXppC7mPHcZ
jEd3OTZR6dcsL4fvSg04AIrc9WYVoyO792IqZQ+zcfbQOYUtDze7+fSRFwRia3qJKLS+zkgH6jmN
NyDVFUGPMFHAESA58yofLQODL8dAtfmvZHyyHcmaIB0bfiIQp+mYGdwvmhKSq7v/iZHJ/utPtegc
mNfPiMpp+ms17EkXepGjIX+0ObPwqLga93lHL57QM3xnNjQUO/ohgSRpNlKYbfYMcS3lNhlHVpV+
TvN+pyPfmJZFBbGrUNRhY4JVkUdk1jUDEYzfkzAGgMZdCEky7rvv/qGzwHLHpZK8xX13OWodRAP1
n8R8kcqxEicCLsJydxFf1tklURg0kFAG+EDiD2YfSJq/A+RLWji+Jy4t98PUzdQ5+TlXWuS3S5kj
cK2Tj8U1W/nuVdkqe9Ox3Tsm0zA1aAPg+81Ik92JmehRUM92WftdIi7vzyORjhcwBIVSHmiHHLYw
Xo3psuuW1mzR3s76s6n23Agtx+EYqrV8IzrTfvC8jZwLzqA3PbRWEJbZNEgd5AB0epFgn7cESnOU
haTQ9s8le1klijQezoagYajSe2I9Qt35H3tJiSX+/kIN2y3ILDsDM1fn7ZT2Hlkz8PQjrEPznJBb
TO69LJaq04TpF+xlHdJpzGPbjpUpmuGFsNm7AF3/LhOOT73NyEOy9uv56zakLxouQmkwEcdtuRlB
PY+p3EiSN2kV+1NLmO4EQ3Bqxkp8YmW++QSs0zSwdpo+Vcgq2edZznaigCM6yNNx9Lsclqo21sfV
qmEYXU0KthcuEa1KFwSn4dwGddobUCE+jtgCRTt3yWnUfEFDtANYWNidFLRmdVWu/pRz3Jvpek6B
uYHQ4y7RzgSuAjKAh/bgbMbRhPfZHse8fHXhQRx2+zSMhTr7cc1rV/6PuOvcGW2bmWZrqCINzzPx
SVSR52E5+Fb0yK/HLrtyfxi2wzGoDEfat0FiR+gTYfIKw9TTOFB2t7RNLO6l0AIEaxXL5kkD5e9h
bT8MQWDlkynRcKgDCldShC03HM/udjEwRd4NONbzFQ8Ow8nxWKLvdG5h5BWsGtAfRMN2vC1vMtiu
80rGcbo6WkRkYgk/tC5gcJigmMSapvJMAjitNmsEJuHQYCRPiugcBSi8mYVRO/f3srFRGBJ/NXU2
CewmDulnqTNw4xWMsVoeKG+s8MJEASRoZAU53wwEA5UEN1RQWXSM9dwH8lUd8XRZFbYX8VYcLNXY
h3fCP9IWZz9LCRmFON1MkVxemCmW7gXq+4pr7vNfeKFTy7YFvAyd7zOM1xci/AZCEFOT3NOJgHEx
jWjrVsUzfFcPGhpfXjeSLrg/GQoqXiMmhstlVbFu7urR/IwUjPOulT6gheF/dcQ1z/suvThkZdWT
6/h51/xyHs42YSFUD8jFMRbtG8heEgF2nnExN4mQHtN6HeI++5tk1hIUW9WFLfpUTlD/be+K0tgj
c5CT19/xM9KSZI4+sGpeC8HFrKHqHJdQYlph8z06DgSzmezVdHmtcZxOQrSGwz0D0xpQBhGhLLgZ
79yVU0DkzbuxJqWpIOrp00pSUykmAS+tw2MId4JAIwMmvccdRmg5KXn1rDEz8g9As8IhCl9/jJwf
Zu5BqbQ/bLhQbqsk/m8/uJjbFewWN6OFha217aMDv2DiZcU34AHr0mrrjzeoaV2bjF5AHg5lcUaU
O6/Vijl50XWb27fEHhQPLsgoJmUzGe9y6q3zfnD9kQo5Qtuf9vjJhUrXV7nHgW+uH6oh2pg+5mg/
TMSSlTfCCnt1rkQH8Leoz7yTKp3QaBmiCji553sSCHHUbq9zBIiEfWlpIOWZDLGF0uRontZdNy/+
bj2XeuIvutHCMSwPvptkmg+qlwDeRPCZF3ZjsSbWOeAafxpuBG+BiGOZNK4VvfgX5zj2T0mBPh9k
e5AQQyM2nHxFeMY8e6q9+7tI+taMuRPrfVTMFlGHOBetc6hcmOA6eduIIzdr4xqSkybvglI2KkcP
BngObzImCaMpeVWYnUTdlIafNMilBlTqFGnfBqPJNU9vQr/OdfS+gRQ3LZStGMc6F1oeHCABML65
g3b7YRhflnL31OtJ3gMIV8fSksfAeeaI+tjnyaBIyyBPcann3dLqrX0Lk5CjnK2u21qZ6jrzAZJg
AROL4HhO4mQW29o6xiE3bxYmuz1Q9x/g7k704ENigmKSCdi49hQjZ7L2CCyTFaoxc51cCAtCatQO
+UUXcEVdNgjXBkjrc2gYtFEg1QLt9077AucpbXS0S2eL3+neeD7/KITzy534Ka2sP2RtAcnB/QP5
3EF37xFthYNf94PikFPYsbUIhcnN74ineiYKzJ6zbY6BzFsK0hLJ15hcUmWnCfi9LVbXQ5QO9vzf
dV6/I9MI+4GfxRN3kE/1V1g2IIZE8hKcoHxBv7rrqY4za3rUhgJS5lP4cxpYQGygouAvpPoH9bbW
N0/XKW8Nrv8yoz6mydRWgucWlNa6EVvjNmLyeSkiCjac6CxyaxmPEgc5o0CUJdX0uc4Vvdj5t88R
5514i5mT1U2hO+1tT3sCxOPJgO/rDKH2YEVDLERmSvuEYt6dVKSEgx5HyxGVdJptMtA5xJtkjCWS
IImeFIvj4or1Osz9pwog6nOlioc1157uIvHJLqsIiuc6krd3539VafYV7RlPwY2bHm/aNFujPUfX
zzDI6eVgfJM0WLDR5BPhEUzGrEEIkk2oovhpDo2eCGCLhvfq3PEiqHgm8IqdLRX8seM6vBG7kjka
zuJXeBipqIAibSYT4cb7swzHq2DA4pnZfNnRiVa3snd+iT8C+dwz8OBgk0qjmPyPVUWzkoNSBa92
11ehrMO8bwA0hZTihLgwnmTevBPvlAzsgTUSEfuLMYezVwyFcjihVtCGzF2VXGYTTbpUzi/8I4hs
Xn/shiDyF8jZGbtiWAkOwD+Q6XV4Dy9haip3uo/l/nR/3LSRT/UVeWUXDLSuoD0BUiGwAXvP1WaX
XYsvAGC9b33UOXZzLGl+FaS67/YhX5r0Yqpn0b08CTb/X7W94JrKOHlVeYLKjlqMEMyezCPDpZ0o
yMGx4JJ6L/QUJSLxLhQHxX5kMYQJvPnkPZTGnCQow10iU2ss0Yqidv2gkxhMmVXktHrgFAe8da//
FsYPSN3MusQtYimZ2+wq7OnwHaX0qq9chYT32o+T3DOlcIn/+NU8G/qpzICZOUQoaJStPj9jWzC2
gSMPbCOUNWe+FrwS5+/Lyf7sPwFu/Tq6vpFKP6gAJDHdq9O/iFYmo+dv2eSZVnQ1ZBfe9Hm0D1Ak
yXsqfat2vytTCQrrLYJAbtje2IrJ1+PBCY6osyO+XlkPHptaMuM7a3tFsJiajqO8BTncu4l+oxt5
2zGl2JhFvaxOBW+ikYmF0KBzqkkCEEsqKhTto99tuFiHGZHPbhxmlPyW/nRpUidzIym2U0H788A0
i+dK3hHrK0jpFFda+b/Hn8tKPvJNzRiR4/jrKds+F9OGdEA9cq9MNm6WnC3sLBrMTya2T3sLchmr
f2L2t/6nx1exNt02rKsvmZJYb7dpuu1zoIbsqCqET4ipyZCge9sgWJ9/8cIiv0AIpbCAeD+wTrq7
JdR60MOtZR8CDZOos736NIO2xgP6Cu/auF9lKze9pVxApx29CHffUuxuzWGe8mXaL6c9hOvT9oGb
bFcB6sYpYor6BxFJjGkdwF8AkG0xWq/KCWtL/VneZPHUbEQFQ7rihMfju7fiXGU6yboOul67B1Wv
wQnH+ERXWga7LcwLT0mKg4hRSvMLpHxI6JEWEpR6fTS/Sg3++MTcrvDVOthBF1uG+2Af+jFySYaR
vBCVBQJoJE/gYgBD3baJFS/i/lToMGYBDjyBPXkaYrGQETmuHLc2s1neZ0QU4Ppf/VLFZd5AEcCy
I4ar6GsnWW6ADgLC4KGgdDvBkCmNlo/2fCatNcEMSDZwh+a1uL20By84FPU2tG6lhdcajK7v/mR9
4dj1KuDXb4LNzdgZrf3JSJsSDaTTh3MHSheIcjU3KobYN9re9PG2r8jMSX2UQwIZNtk4a0oOHpKt
RQiHCdGOxnY5R87EtlgX0Q1wgkXFYyO30VZT6AQBCIbPBFOVpGh+yYcd3pnzQ06nOhcdKV6Ga01B
DvIavoInfwVH/zYtXapnZBttl8mklCV94gn7P6fZBQYRDBs/e02eGGnunoitMqF5ekoGOZAwbzkp
ql1taXV4gofDyQuSf6edF+mQnpx3CIirBLdM+z5oevOAciy59t3TgxjuURk7LgjGPQWdRKmF6T22
ffrFMD8jeFW8AWpuxmn1fEEynDGtIK2Gv3t5l94rbay0FJXObYuk4duZFvKqwZosxqLq1PvO7vo4
OpXX5yKtpw2+AI86eijWEQ5/z9qRlF4USxAyAPEb+h0KIkCdEQAYXdW6ywwWMUYv3gsl/B3QIHSQ
G9VFeLsyhcqcCfas03SXQP/q/764RMTieEfo5a6LNB1QRuw763cANCamNWTenqBvmaH7KYFzjcpP
7u7wt/AtMwQ73KAgpw+FFE4e1mp1+K9W1/Lb94o0mxIfroKknlz9zq5xwHehEtZz3M++yox+EXWI
ytfSIzOIEMN/jkML7KyuK9t084CcMq6QOJYvx+dybU0akwhZ4e1zMgBCe5SuCgjxd6rgOOlVRsKf
c8O1NCpJjU/fV/Zd3nO2kmnfuZ45PDdJLonx03+d+vvvtuSQ4ygYPPBmRJwo8DNcypgAzvz+1Geo
7/rXizk2+wBkyQAl/3fIqUs3FNKcHH97jg/UnrLlGRBLOszAcoRw2MNADyRxv5PZXgL+bnIq1fXV
ynAZCrZ7I/1bb63nufXEnWCpjXKwEdjMD1Nlq+8jhRY0aCHMAfHiVOkVRHp+WT+qUqHjZ8WFDNX+
OAetK9DGijbWWjpN3nOrxndzEDlNgmgj1DQISolI2gLqBaW9xgvhsTacIKWcJE6LC2gvk2SmblU5
g/cOikO7siX6r8Nx28saDJ0UjR01W2JJaDBLkkuscf0vy6drB4pPcjyB6Xly+gk4y7jFWm953qOr
k7qIQ+Ia0rHvm7RTER3jRWZrZGpO4K7KwmejE6zumepHJQv9MjCIxm541EMSMQnFC2c9QDpFMTtA
RkGtNUlvgV31uIWclIxN08hWM3tcpUGffL9klbT6k9FysBqRTBQPh+3zpyCKVSVBL+REb9d7o1cR
+qiMLaPFdu8gjywJu019QzXDl3+vYEp8Ny7Py+5DYkOTt2wMiLCZQ9kDhvVypY9eNUXnhz7tO5iB
TdO55fuOcnMLQrvT/pYNlYXswuY+/qzZVi5OUkRWvE+cfoZMGmy92VWyzLG9mYFen8IgM49NFrnq
+E8AMzOsTxSqdtqo8k29bwKgOjmSXKAfRItyhCaHdORWe03Z1T2hlakmQLY0CHhYLw0Ypf8QrO4k
WxCcs7rf833JGUjl/dOaGHsuImrGxQoJuxlelrCsVewyEzoUgwpSo/EGJEuhXgfHyDwSwDCk62Y6
wmNqdtEMNvJF303r0lIXYUiJ1nt33CLWqZ03Ev3z5f08JO8nrt8OMQj0IGr4/FOSB4ApHNJ7VQaI
EOljZ8qh4lvLB4SJmWpH51eS0q4bfDyQV6y7otaYMRqhlZnFkgxJQa/A9BENf9Uf7137oX009Bwu
fZyTAbFWb/suViIMDijAufOdAyEIpCKKFYrTy70Nw/kf+OvfGYGu2br6B7iGzJ9ziQKFZpSweXRw
2FE9A1ZzCWaltLy+xEPJYH80VKX8aujn+yCl8gwob0Dtdt30gWhx0+YS/rvs0z+F10X46BQhU0sX
DGN3MFmdonAbvL2/R2OthBNt2RC+qyj5zG2l3tg96a+4KcHxVkm52hLFZdSm8CfvWEMv0XYDaj+x
pNYLADtniM/YcaYdYgzuOIorlgcALdtJ2gePfa3Gp85e8BvAd9HSeQtsJg/ugjusmOxe4FrsWvy7
MAQe4qByEBGG3jejgQEsdwPblbXm2FumGjLpDLDqxxEfpqqTRuI23H5Om5jmxkK6ghoeUcDJT/EY
tb5TGGDq1VtkJZef2BQnGG0bKKbez8Mg6FG2oRIbWkGhkSZBXbD0/iqn1CuwZnuAhu4Z3Uim4N4/
nlSo/HKj2WAp1eE/79LCSBRa2kSnfGJ4WXGXFUQ/vCcVJiq9r2B85FrIN/DujRsYC2nC7Ux9JjS3
mdKeBUmUuI2ztII0s2odlORAoWNRTHOugrXOygMNKMTdNIipSHIhijB3LkWM8enq80kjO9qdrrIv
x22/xoTJnEK5Jhf8DcWa58kjuwMOfYf7OzbgmczdyaTLS7+eU23RHWonyilDDuZPF1fGRz8NklII
wagk6eP6pQcoqDXKYCMwPyjTlYA/iMqCvedpDMLuUDDyE77WmBx66OC6tOlEtmucl3F4vuNFS62D
H8LiqSoA8wRdZgIY/cNdltnPudT18SIS4bGaBB8hSkBdOBGyNd6fbWgkesqjwrEka8BxuC9bTdI6
R0K0auHIfzcT/XdI1nDJtMY0Kayy+lmVdM6Xg4Zl2SnbA5ot9fKCNJci3I55kqsyogDqXGGWulnQ
uFmrUHqI5HWlsCDPFH0uCux5xIAYQMOEK6Ek6mQ4rZJ05vNkQeyNc7FWjX7keH2sMU48LUOhO8Q0
siLd0gPI9VtPF2ZxDxUnY16toXwaDE4Ah4m8e7ydsOALoUQ2J90sDsIabPATfzB4D3grc7Z2x1pX
HXttV2D4DLNwp9eV5JHjpYRSwm6g+lkCoo+dxVqaR2Du9u8ZUAlZkCGXkxcjLNQ6eh106zXBRPmd
el+a6Qez4cAHFPezrv51pZJUqRvrPjMFNGRl+j0TcqS4/sw5E5V1/2uFtC7AD0cDythEx+iOBzHd
u2H9FPiHnJ/I2VZRHoz7qM7l6hm5EqAPfT27iNEMu3JbqbgqBlnP3CKBmy9nrQjnp+qTU3QMaoUx
soD4rlng5yoPyRKJduBpTnfHx3bKKkQZ57Ad4F20l18Imo/EWGhdogtTrNkW6sByxa7GkiHIYpF0
WYkmmTdSS5fa9kcB53PTdH+PeyS6Rao4Zf6vVd5SBW1jslV/X6FWWa+PRZ2GtQ7OzMck1hwBXyan
lPKzmboh6GLvQgAUQLg0oM+NQJNTuUqHGuxB8+LapTNEM0YUQD0Z01g+AOgrDctVFPg8jUAqV7Zl
0p/teAlaXkq/Vt5zP6t73JwmqEi0mkFcFOniiRzDPouUaEWsb5ioQ6BK5phVegyCwGg8NSo5/SNh
L+MRO3r+QDrbPFQ3H2TbpLAUa0HfNTChmkRYK/kQmMlgMz9FNIEQHnGl3+P5S+xmM7sb09ATfBko
ICx/sSoF/MFNdxxnbq9mUUihoW0UMCxjHQSof3331B/jXfJM0ghY4HbXH8yOS3uKFL4iWQc68f7j
bI3TDicpcrE+HGBIHs9671OHh8jpOEdpYROjEytnvs5nJ3WHK4RTrA/vN/wlyuNmAdeWo2mSw6tP
X61CUzdwCoOlDxMaoze3C+6oCJcfIjQsN5t6m97Awc3hWkSO3k84FaEjXk50Yb5Qavvt7nNuwpEP
2v13hN5DBvdRmBwMF1zKM/S7me49EvP9SuoNZCCkwwe4QdtWw3glHBWkoiXy9PZKkkKMbshN5gzx
o4Xdlra/lYFbTcq1LzTIN3twgpRQaAujvOpc6VWxHaTASbVzII4QJrLNuKFmYVAExvQgwAN05Ece
XZZNHpw9Ac0RSbkfAbjYk9226pjzljOP1twgyGax2fNrla3fyDBWmIm4rhUMR/HO/NMRkGBCmHZH
YNJT9knhYOTpVtsEWn05Rc8UDVlZCRRdX7P6OzLTDbwboJMSEVGu500toVLPuQyoA9Q6MDw/lpBf
IFTTRa7O1jMAq+7s1fXLhGomtc/dMddFuAlC/0wuWXx95fF5zqT0Oz65olsGbYEEPHJaYC4JWEPb
fEIjuihtuer9k8XvKutsAlxcJE9eTAwS7TMjuQ/mXVslBWGJUoF7YxZnizoAGU/ayzCDazKRlYzs
Bhf24jVlzOnqwVM7EgHKwlL+1MC5TCO2/3JqSN56Z4Ze4NixrQpcnHTsbV9CpLrcggWxvQGcwm3U
rB4bDNZ78vDgrpNVohtBqObBes8D/YkjPPkl79RBckEU9Z7rUzsNUf8bKs9kbL+qABQqbDCVGkhH
6BHA0jDJxOvUyJAd8UaADgcU2vDlUcZigT4MkwLFoJb588T+ktts9Cd3K7PvpV6my7AOGUQjqdoR
SFPni5ISzipi4l5mkP4aRRD/1PizqPDepbuIZvdvRbOkih4TN8bVZ439V29mC0uB2eSv0FkO9uzU
aUCo2bIozNZw9O3UNaAJzjLm96Z8nvr2Pbk/f2js2mn1Qrgp+avAM3raB/wQRnssr22iUvhkuK6L
Q36jA9ScShcsIA5kDIr5dwGLNcw9hvwa8uZvEipegJOVulpGCqV+vygOJE4JvS+HtouCKyOu5dyD
zsdjcbjMAy3RE1yNutZv7SEk6Ze8B9pmPr4XEWZrR1KDuTKbByE2P0jKbJbx2/wdfSnBdPuE0STO
zPIQuFN512NvgRmT/c/pg7yjv06JOAAzQ85qLV7PZ5K/suEzzjU8ImFKu0HKElke+NsFUUsKst1p
dP3ZSENGnFPWlTxPtBlbbiPCeEUw0HEefu9jHUAknGgWPURkG3IHYz+Fr4xqicyd9adjCfrO/rn4
W0DJrYvKYeCV+Xhvp4yS0Asw4R/vs+msiMU1VBv/5mOap8lYqL/uImI+WYyK62cDHX1dX9mQLkJH
G/pFMLhlyCuuREZeJCKHllKysub2r5pnk1FHZiiV7jz3a73sXplnkDf/a57B72Qz44NcXXdiJ5JP
qUKmoVq520IpyGcwhHGTAbgOYp/vdbKmFiYdBCNwzjXH/x5MOgyjH8Qi9CQQ51n4t9lGqqygQeqQ
WADLjfY0ZXfHA1+4vkCSlu9Azc/Pz3i+mCFIDeykJbjKeKhEc6dVZ3FkRUJsboJYj7LEsyxQC8hk
c3RTiHfwYslBHw0FaQUi/Mbz3hZ21r9Rk7uFLkKx9No47sUIwCfEVBdms3SmDQZ2wZ22dMyJXaEQ
wtpn33w6fNGNI4PYGlA84jUTQJrqoIMh/DLBmr0JrL3i3cmXtpU75jC0wG/JekVX9qP+2Mb8HG5S
GfWWftCjS7fTw4PG4DXiK/Ypx5XM1N060tJ0lU+yWbhzM6shih7joS+0uQDYNE6fVfwymNaHvJo7
i7lpS3JERt7YNG5IyffJgTg+vz3PTdKxDnoEy/6p+04RNjXeaws1iYcrJGEociM9RWO0WmXUP70u
fymoim/PalxrTtbFxi7H51uHtvfP+aHygiIiUyJWjSR5Sib4fNl7QBaKleLJt0PK52S+uVcmBUSj
hpOj2kJX2+57ZzR2tkdD4m327Z+0kl9ALTxRrEoP/k5uPAjyUkb07WIrHB9wYxo01tgcqn7ToP3w
a9A3fOye3PEMOvRbD3C2KfUHc41T3FzzPMVlLHTnzx6Nwq3r7AZARpPgsMbRSA7v01y/fUyhegvk
3uTr4FrwSPG7Sia6EhVR5lumxUabT5zBz940EHIz07QRSttLW2RP3eJOkpNKgwJSQFqPbl02ItkR
oBn4kq/6rCeG9k2/Qp56duc4YdThzcQxUaNa4XbIrlwU9sPFY3LSknlzx3NeyOgYISpGmZdHzomU
SIlSXt9E0jc6f3M5fitDCDCIFvlZ+gvGFS3Qr0SlqcZiTv9azWdn3UxWeiFxGCCSfwdWiY7erw+T
gQnD+vQkwLFZH7TWbNmuyHcF58OolmYaGjZsRtTn29eJllBo56t9JL+O4ugA+dPb9cTTiGDdUy7l
TSSt0kBr3DKc+BzBLlDdq5R6QuMcbjB9/5h0g+WPqKogHwph5E9Qo1J5gqtqMxE8iKsdu815qvzz
P4duMWY3QuY63W3VKawrxTpq/2vIEV2nmd8NzcDKw/1x2Cj+GZ8eouwMepwdmPZ62benWP2YdaET
xoJ+4P/LYJYY5kIJadcfdHISJinXMZggI13UT2BBesHmTc1KlDDiHDX22HviucDDi4jzfxxCvgfd
ELx6ZfmunudOwQyR0vnTcieF8yj1qdEMCS/NrLnLTrf4OoyzNcXLbY2RSbjY1wnWylnd9nIm/tLb
5uG+POPr4M5Hu1VlIu7qijl/LmMfBiSWq4vUEnD/8ewMtlpcMf0Mw1mD9v/7mgsJ62/u6d0/m7ND
uEm6fFmjfUdUPm2YLCA70AeyPkp3li9H0rf0RO8Bs5En6n3Q012sOVb74DcStTABS5F8eZ5o14W0
mP3j5FVfGblTKoYvTjJzzyNHjxrXEY6N1yh8GWN5UruawAgRsMVRn6DT1M/5krkkT7oEb5MMdNYq
663/+EXoukDMoFvEfhKJZOPsiNVMlqnvm/qzv1gSpcTWbXR1ENtxBe8RYyrrUX2RyR4UDAyKaU+w
w4sVpeVhYO/VCvpixEe2BUTQ37LKd23L64WB20Bb76Ishv4kQd0e3z+EdN5guEuLaQqlIeItcO9t
92dyBXIq/VEVAAsyJYZlAahOcq+6vUprcEwFAXl2+cPiP+RY5Yf6vFPmCoc0un5J0vEgNn/Elb2h
3Jr6IIcHLMGEba36NS79Hth0bYN/OkTR89lK+3ZaTVDGjRkjqx60KA5ToFB+VNb7rYwQn/sZzkZ+
k0EcOaoU8QOnKz8cTI4tNnAwCnVK4cuSsL85zUijoK6aJSnktKY+rJL8c6Ti7I2I7U/a0CsG0QIu
jaSqqmhI4td819XTVSEVKbMkhq7YCkdUULKr+TAXFgqNBNwGAyjy+w/Mgk2ziiyMMBv2WpCt0E7j
F1QlXRLqd4UVJ/3k4brsS/qMA7aibVXup+23EMKSbwADiESvWXnLJIOJxJuK+ZGLHn9S5dAS0Zy7
3SymsgUI8pLJ8WJ4NeVfnYChBKAtoOiHArRsaYRL1LMmjEsrSpbMopf3n2pstCbOWBBcxVFfp/Jx
kbeza6hYJ+bg6qygBeblzcvL1F7W0ilcXRPZcTkAKwsbmzaQ5UJWSCFvmMwhyFroqCHUvsO0PimN
mO9qM8sNHnoEj0OLWcrXu5JybpqB+JWTKCIJEo4kI3SW5ugkJG7CM/ykSjs9cjQ1fHCSvbULfzBB
9c90Q6lIFKPa/ugtuHyD5eCmp9ePQsP35QY451ZQ8UITIYoKXkcHzls+khtfbJTo071KLEGTe+pD
qk8jlbgdcr+DQ4ebvJ/up25Yrj9JC4NAw+kaN/VU8NAq/ogwmeaiWdSiooQj6bZt8t22vi+GxEkI
eYzdX7MASX9FNyVfY0AoDpG2IiRkZ3kD3d7clv8z/1Q7Bbts5Nas5V9O9TdaiU4BvvwgnGs5eI8d
kQGwkQDWUdUiXB2t5bfVLF39vkcTkbrhjdRWpEYOojqSq21CemfHPfZevUlBLZfPtbvE5jKFWcCK
PxivZ8YtiZRGdj5EKbuIyPKbEfu4ti6EDxYEKJ+hsrhQlAcamYSVoSkwejK9AC6zxEFt2LmarKXA
NEt1/1ZzYO2i4h0LkxxVCULv9o4JjBv+BMZLaGG7fPctJzIOL//qSzyjiZiMYwgm7OK5V4n9gGVS
ggVdAVpZ7x1xbSwtlA2Q9FAryjEcmJaPHiqjhcB+EpdAaEs=

`pragma protect end_protected
endmodule