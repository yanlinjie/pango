version https://git-lfs.github.com/spec/v1
oid sha256:d4a3139308e557cdad84712b6fa0ef6a27e267359e0b635c5f669823c84a9209
size 886
