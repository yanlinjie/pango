version https://git-lfs.github.com/spec/v1
oid sha256:f0962a0e6983bc4e47b9c27e7d0e94a7d5e3c977c84ba0647ad622f45176b4b8
size 1163
