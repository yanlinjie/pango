version https://git-lfs.github.com/spec/v1
oid sha256:58d41f3cdfb80dcabb8ec1637779c1aa615c7152afcd2fc75113415cf471f518
size 582
