version https://git-lfs.github.com/spec/v1
oid sha256:e93d207748abaff5406e6243d34c6b1696dc1f6a1716cca7f9a256146376ab6e
size 86711
