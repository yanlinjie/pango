version https://git-lfs.github.com/spec/v1
oid sha256:301584d05c947d0186153d94274781ea8b86dd91946b0365150f46907228d1bf
size 1269
