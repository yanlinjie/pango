version https://git-lfs.github.com/spec/v1
oid sha256:e27f51d7db65076782f921f9dea0e20ac26ae2a5295f69d02d6ec7ee8d82fa3b
size 1069
