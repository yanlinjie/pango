version https://git-lfs.github.com/spec/v1
oid sha256:ad9ccc2beb5a98aa13db623772b7721eb0d5c4af6433cd0ff5b38d00c4eaa02e
size 1263
