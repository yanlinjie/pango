version https://git-lfs.github.com/spec/v1
oid sha256:1a362e165229c239796b3c1d7f1e99433d461620b04391fb7af0da4d9df216e1
size 1269
