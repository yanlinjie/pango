
//////////////////////////////////////////////////////////////////////////////
//
// Copyright (c) 2020 PANGO MICROSYSTEMS, INC
// ALL RIGHTS RESERVED.
//
// THE SOURCE CODE CONTAINED HEREIN IS PROPRIETARY TO PANGO MICROSYSTEMS, INC.
// IT SHALL NOT BE REPRODUCED OR DISCLOSED IN WHOLE OR IN PART OR USED BY
// PARTIES WITHOUT WRITTEN AUTHORIZATION FROM THE OWNER.
//
//////////////////////////////////////////////////////////////////////////////
//
//  REVISION:
//  15/06/2020  mm/dd/yy - Initial version,                                                   
///////////////////////////////////////////////////////////////////////////////
`timescale 1ns/100fs 

module ipml_hsst_hsst_test_wrapper_v1_4 (
    input                P_REFCLKP_0,
    input                P_REFCLKN_0,
    input                P_REFCLKP_1,       
    input                P_REFCLKN_1,            
    input                P_RX_SDP0,     
    input                P_RX_SDN0,        
    output               P_TX_SDP0,
    output               P_TX_SDN0,
    input                P_RX_SDP1,                                
    input                P_RX_SDN1,        
    output               P_TX_SDP1,
    output               P_TX_SDN1,        
    input                P_RX_SDP2,                                
    input                P_RX_SDN2,        
    output               P_TX_SDP2,
    output               P_TX_SDN2,  
    input                P_RX_SDP3,                                
    input                P_RX_SDN3,        
    output               P_TX_SDP3,
    output               P_TX_SDN3,  
    //if with user logic
    input                P_RX0_CLK_FR_CORE,       
    input                P_RX1_CLK_FR_CORE,         
    input                P_RX2_CLK_FR_CORE,         
    input                P_RX3_CLK_FR_CORE, 
    input                P_RX0_CLK2_FR_CORE,
    input                P_RX1_CLK2_FR_CORE,
    input                P_RX2_CLK2_FR_CORE,
    input                P_RX3_CLK2_FR_CORE,        
    input                P_TX0_CLK_FR_CORE,       
    input                P_TX1_CLK_FR_CORE,         
    input                P_TX2_CLK_FR_CORE,         
    input                P_TX3_CLK_FR_CORE,
    input                P_TX0_CLK2_FR_CORE,
    input                P_TX1_CLK2_FR_CORE,
    input                P_TX2_CLK2_FR_CORE,
    input                P_TX3_CLK2_FR_CORE, 
    input                P_HSST_RST,
    input                P_PCS_RX_RST_0,
    input                P_PCS_RX_RST_1,        
    input                P_PCS_RX_RST_2,
    input                P_PCS_RX_RST_3,        
    input                P_PCS_TX_RST_0,
    input                P_PCS_TX_RST_1,        
    input                P_PCS_TX_RST_2,        
    input                P_PCS_TX_RST_3,
    input                P_PCS_CB_RST_0,
    input                P_PCS_CB_RST_1,
    input                P_PCS_CB_RST_2,
    input                P_PCS_CB_RST_3,
    input                P_RXGEAR_SLIP_0,
    input                P_RXGEAR_SLIP_1,
    input                P_RXGEAR_SLIP_2,
    input                P_RXGEAR_SLIP_3,
    input                P_CFG_CLK,
    input                P_CFG_RST,
    input                P_CFG_PSEL,
    input                P_CFG_ENABLE,
    input                P_CFG_WRITE,
    input    [15:0]      P_CFG_ADDR,
    input    [7:0]       P_CFG_WDATA,
    input    [45:0]      P_TDATA_0,
    input    [45:0]      P_TDATA_1,
    input    [45:0]      P_TDATA_2,
    input    [45:0]      P_TDATA_3,
    input    [3:0]       P_PCS_WORD_ALIGN_EN,
    input    [3:0]       P_RX_POLARITY_INVERT,
    input    [3:0]       P_PCS_MCB_EXT_EN,
    input    [3:0]       P_PCS_NEAREND_LOOP,
    input    [3:0]       P_PCS_FAREND_LOOP,
    input    [3:0]       P_PMA_NEAREND_PLOOP,
    input    [3:0]       P_PMA_NEAREND_SLOOP,
    input    [3:0]       P_PMA_FAREND_PLOOP,
    output               P_CFG_READY,
    output   [7:0]       P_CFG_RDATA,
    output               P_CFG_INT,
    output   [3:0]       P_PCS_RX_MCB_STATUS,
    output   [3:0]       P_PCS_LSM_SYNCED,
    output   [46:0]      P_RDATA_0,
    output   [46:0]      P_RDATA_1,
    output   [46:0]      P_RDATA_2,
    output   [46:0]      P_RDATA_3,
    output   [3:0]       P_RCLK2FABRIC,
    output   [3:0]       P_TCLK2FABRIC,
    output               P_REFCK2CORE_0,
    input                P_PLL_REF_CLK_0,
    input                P_PLL_RST_0,
    input                P_PLLPOWERDOWN_0,
    output               P_PLL_READY_0,
    input                P_LANE_SYNC_0,
    input                P_LANE_SYNC_EN_0,
    input                P_RATE_CHANGE_TCLK_ON_0,
    output               P_REFCK2CORE_1,
    input                P_PLL_REF_CLK_1,
    input                P_PLL_RST_1,
    input                P_PLLPOWERDOWN_1,
    output               P_PLL_READY_1,
    input                P_LANE_SYNC_1,
    input                P_LANE_SYNC_EN_1,
    input                P_RATE_CHANGE_TCLK_ON_1,
    //Lanes
    input                P_LANE_PD_0,
    input                P_LANE_RST_0,
    input                P_RX_LANE_PD_0,
    input                P_RX_PMA_RST_0,
    output               P_RX_SIGDET_STATUS_0,
    output               P_RX_SATA_COMINIT_0,
    output               P_RX_SATA_COMWAKE_0,
    output               P_RX_READY_0,
    input    [1:0]       P_TX_DEEMP_0,
    input                P_TX_BEACON_EN_0,
    input                P_TX_SWING_0,
    input                P_TX_RXDET_REQ_0,
    input    [2:0]       P_TX_RATE_0,
    input    [2:0]       P_TX_MARGIN_0,
    output               P_TX_RXDET_STATUS_0,
    input                P_TX_PMA_RST_0,
    input                P_TX_LANE_PD_0,
    input    [2:0]       P_RX_RATE_0,
    input                P_RX_HIGHZ_0,
    input                P_LANE_PD_1,
    input                P_LANE_RST_1,
    input                P_RX_LANE_PD_1,
    input                P_RX_PMA_RST_1,
    output               P_RX_SIGDET_STATUS_1,
    output               P_RX_SATA_COMINIT_1,
    output               P_RX_SATA_COMWAKE_1,
    output               P_RX_READY_1,
    input    [1:0]       P_TX_DEEMP_1,
    input                P_TX_BEACON_EN_1,
    input                P_TX_SWING_1,
    input                P_TX_RXDET_REQ_1,
    input    [2:0]       P_TX_RATE_1,
    input    [2:0]       P_TX_MARGIN_1,
    output               P_TX_RXDET_STATUS_1,
    input                P_TX_PMA_RST_1,
    input                P_TX_LANE_PD_1,
    input    [2:0]       P_RX_RATE_1,
    input                P_RX_HIGHZ_1,
    input                P_LANE_PD_2,
    input                P_LANE_RST_2,
    input                P_RX_LANE_PD_2,
    input                P_RX_PMA_RST_2,
    output               P_RX_SIGDET_STATUS_2,
    output               P_RX_SATA_COMINIT_2,
    output               P_RX_SATA_COMWAKE_2,
    output               P_RX_READY_2,
    input    [1:0]       P_TX_DEEMP_2,
    input                P_TX_BEACON_EN_2,
    input                P_TX_SWING_2,
    input                P_TX_RXDET_REQ_2,
    input    [2:0]       P_TX_RATE_2,
    input    [2:0]       P_TX_MARGIN_2,
    output               P_TX_RXDET_STATUS_2,
    input                P_TX_PMA_RST_2,
    input                P_TX_LANE_PD_2,
    input    [2:0]       P_RX_RATE_2,
    input                P_RX_HIGHZ_2,
    input                P_LANE_PD_3,
    input                P_LANE_RST_3,
    input                P_RX_LANE_PD_3,
    input                P_RX_PMA_RST_3,
    output               P_RX_SIGDET_STATUS_3,
    output               P_RX_SATA_COMINIT_3,
    output               P_RX_SATA_COMWAKE_3,
    output               P_RX_READY_3,
    input    [1:0]       P_TX_DEEMP_3,
    input                P_TX_BEACON_EN_3,
    input                P_TX_SWING_3,
    input                P_TX_RXDET_REQ_3,
    input    [2:0]       P_TX_RATE_3,
    input    [2:0]       P_TX_MARGIN_3,
    output               P_TX_RXDET_STATUS_3,
    input                P_TX_PMA_RST_3,
    input                P_TX_LANE_PD_3,
    input    [2:0]       P_RX_RATE_3,
    input                P_RX_HIGHZ_3 
);

wire                P_PLL_TEST_0            ;
wire                P_PLL_TEST_1            ;
wire    [5:0]       P_RESCAL_I_CODE_O       ;
wire    [3:0]       P_CA_ALIGN_RX           ;   
wire    [3:0]       P_CA_ALIGN_TX           ;   
wire                P_RX_LS_DATA_0          ;   
wire    [19:0]      P_TEST_STATUS_0         ;   
wire                P_RX_LS_DATA_1          ;   
wire    [19:0]      P_TEST_STATUS_1         ;   
wire                P_RX_LS_DATA_2          ;   
wire    [19:0]      P_TEST_STATUS_2         ;   
wire                P_RX_LS_DATA_3          ;   
wire    [19:0]      P_TEST_STATUS_3         ;   
wire                P_RESCAL_RST_I          = 1'b0;       
wire    [5:0]       P_RESCAL_I_CODE_I       = 6'b101110;
wire    [3:0]       P_CEB_ADETECT_EN        = 4'b1111;
wire                P_CTLE_ADP_RST_0        = 1'b0;
wire                P_TX_LS_DATA_0          = 1'b0;
wire    [2:0]       P_TX_BUSWIDTH_0         = 3'b0;
wire    [2:0]       P_RX_BUSWIDTH_0         = 3'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_RX0   = 8'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_TX0   = 8'b0;
wire                P_CIM_DYN_DLY_SEL_RX0   = 1'b0;
wire                P_CIM_DYN_DLY_SEL_TX0   = 1'b0;
wire                P_CIM_START_ALIGN_RX0   = 1'b0;
wire                P_CIM_START_ALIGN_TX0   = 1'b0;
wire                P_CTLE_ADP_RST_1        = 1'b0;
wire                P_TX_LS_DATA_1          = 1'b0;
wire    [2:0]       P_TX_BUSWIDTH_1         = 3'b0;
wire    [2:0]       P_RX_BUSWIDTH_1         = 3'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_RX1   = 8'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_TX1   = 8'b0;
wire                P_CIM_DYN_DLY_SEL_RX1   = 1'b0;
wire                P_CIM_DYN_DLY_SEL_TX1   = 1'b0;
wire                P_CIM_START_ALIGN_RX1   = 1'b0;
wire                P_CIM_START_ALIGN_TX1   = 1'b0;
wire                P_CTLE_ADP_RST_2        = 1'b0;
wire                P_TX_LS_DATA_2          = 1'b0;
wire    [2:0]       P_TX_BUSWIDTH_2         = 3'b0;
wire    [2:0]       P_RX_BUSWIDTH_2         = 3'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_RX2   = 8'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_TX2   = 8'b0;
wire                P_CIM_DYN_DLY_SEL_RX2   = 1'b0;
wire                P_CIM_DYN_DLY_SEL_TX2   = 1'b0;
wire                P_CIM_START_ALIGN_RX2   = 1'b0;
wire                P_CIM_START_ALIGN_TX2   = 1'b0;
wire                P_CTLE_ADP_RST_3        = 1'b0;
wire                P_TX_LS_DATA_3          = 1'b0;
wire    [2:0]       P_TX_BUSWIDTH_3         = 3'b0;
wire    [2:0]       P_RX_BUSWIDTH_3         = 3'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_RX3   = 8'b0;
wire    [7:0]       P_CIM_CLK_ALIGNER_TX3   = 8'b0;
wire                P_CIM_DYN_DLY_SEL_RX3   = 1'b0;
wire                P_CIM_DYN_DLY_SEL_TX3   = 1'b0;
wire                P_CIM_START_ALIGN_RX3   = 1'b0;
wire                P_CIM_START_ALIGN_TX3   = 1'b0;


GTP_HSST_E2
#(  
    .PCS_CH0_BYPASS_WORD_ALIGN                ("TRUE"                        ), 
    .PCS_CH0_BYPASS_DENC                      ("TRUE"                        ), 
    .PCS_CH0_BYPASS_BONDING                   ("TRUE"                        ), 
    .PCS_CH0_BYPASS_CTC                       ("TRUE"                        ), 
    .PCS_CH0_BYPASS_GEAR                      ("FALSE"                       ), 
    .PCS_CH0_BYPASS_BRIDGE                    ("FALSE"                       ), 
    .PCS_CH0_BYPASS_BRIDGE_FIFO               ("FALSE"                       ), 
    .PCS_CH0_DATA_MODE                        ("X16"                         ), 
    .PCS_CH0_RX_POLARITY_INV                  ("DELAY"                       ),    
    .PCS_CH0_ALIGN_MODE                       ("1GB"                         ), 
    .PCS_CH0_SAMP_16B                         ("X16"                         ), 
    .PCS_CH0_FARLP_PWR_REDUCTION              ("FALSE"                       ),    
    .PCS_CH0_COMMA_REG0                       (10'b0000000000                ), 
    .PCS_CH0_COMMA_MASK                       (10'b0                         ), 
    .PCS_CH0_CEB_MODE                         ("10GB"                        ), 
    .PCS_CH0_CTC_MODE                         ("1SKIP"                       ), 
    .PCS_CH0_A_REG                            (8'b01111100                   ), 
    .PCS_CH0_GE_AUTO_EN                       ("FALSE"                       ), 
    .PCS_CH0_SKIP_REG0                        (10'b0                         ), 
    .PCS_CH0_SKIP_REG1                        (10'b0                         ), 
    .PCS_CH0_SKIP_REG2                        (10'b0                         ), 
    .PCS_CH0_SKIP_REG3                        (10'b0                         ), 
    .PCS_CH0_DEC_DUAL                         ("FALSE"                       ), 
    .PCS_CH0_SPLIT                            ("FALSE"                       ), 
    .PCS_CH0_FIFOFLAG_CTC                     ("FALSE"                       ),      
    .PCS_CH0_COMMA_DET_MODE                   ("COMMA_PATTERN"               ), 
    .PCS_CH0_ERRDETECT_SILENCE                ("TRUE"                        ),    
    .PCS_CH0_PMA_RCLK_POLINV                  ("PMA_RCLK"                    ),      
    .PCS_CH0_PCS_RCLK_SEL                     ("PMA_RCLK"                    ), 
    .PCS_CH0_CB_RCLK_SEL                      ("PMA_RCLK"                    ), 
    .PCS_CH0_AFTER_CTC_RCLK_SEL               ("PMA_RCLK"                    ), 
    .PCS_CH0_RCLK_POLINV                      ("RCLK"                        ),              
    .PCS_CH0_BRIDGE_RCLK_SEL                  ("PMA_RCLK"                    ),      
    .PCS_CH0_PCS_RCLK_EN                      ("FALSE"                       ), 
    .PCS_CH0_CB_RCLK_EN                       ("FALSE"                       ), 
    .PCS_CH0_AFTER_CTC_RCLK_EN                ("FALSE"                       ), 
    .PCS_CH0_AFTER_CTC_RCLK_EN_GB             ("TRUE"                        ), 
    .PCS_CH0_AFTER_CTC_RCLK_SEL_1             ("PMA_RCLK"                    ), 
    .PCS_CH0_PCS_RX_RSTN                      ("TRUE"                        ),       
    .PCS_CH0_SLAVE                            ("MASTER"                      ), 
    .PCS_CH0_PCIE_SLAVE                       ("MASTER"                      ), 
    .PCS_CH0_RX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH0_RX_BRIDGE_CLK_POLINV             ("RX_BRIDGE_CLK"               ),   
    .PCS_CH0_AFTER_CTC_RCLK_EN_GB_1           ("TRUE"                        ), 
    .PCS_CH0_PCS_CB_RSTN                      ("TRUE"                        ),                 
    .PCS_CH0_TX_BRIDGE_GEAR_SEL               ("FALSE"                       ), 
    .PCS_CH0_TX_BYPASS_BRIDGE_UINT            ("FALSE"                       ), 
    .PCS_CH0_TX_BYPASS_BRIDGE_FIFO            ("FALSE"                       ), 
    .PCS_CH0_TX_BYPASS_GEAR                   ("FALSE"                       ), 
    .PCS_CH0_TX_BYPASS_ENC                    ("TRUE"                        ), 
    .PCS_CH0_TX_BYPASS_BIT_SLIP               ("TRUE"                        ),          
    .PCS_CH0_TX_GEAR_SPLIT                    ("TRUE"                        ), 
    .PCS_CH0_TX_DRIVE_REG_MODE                ("NO_CHANGE"                   ),          
    .PCS_CH0_TX_BIT_SLIP_CYCLES               (0                             ),         
    .PCS_CH0_INT_TX_MASK_0                    ("FALSE"                       ),              
    .PCS_CH0_INT_TX_MASK_1                    ("FALSE"                       ),              
    .PCS_CH0_INT_TX_MASK_2                    ("FALSE"                       ),              
    .PCS_CH0_INT_TX_CLR_0                     ("FALSE"                       ),               
    .PCS_CH0_INT_TX_CLR_1                     ("FALSE"                       ),               
    .PCS_CH0_INT_TX_CLR_2                     ("FALSE"                       ),               
    .PCS_CH0_TX_PMA_TCLK_POLINV               ("PMA_TCLK"                    ),             
    .PCS_CH0_TX_PCS_CLK_EN_SEL                ("TRUE"                        ), 
    .PCS_CH0_TX_BRIDGE_TCLK_SEL               ("TCLK"                        ), 
    .PCS_CH0_TX_TCLK_POLINV                   ("TCLK"                        ),                 
    .PCS_CH0_TX_PCS_TCLK_SEL                  ("PMA_TCLK"                    ), 
    .PCS_CH0_TX_PCS_TX_RSTN                   ("TRUE"                        ),                 
    .PCS_CH0_TX_SLAVE                         ("MASTER"                      ), 
    .PCS_CH0_TX_GEAR_TCLK_EN_SEL              ("FALSE"                       ), 
    .PCS_CH0_DATA_WIDTH_MODE                  ("X16"                         ), 
    .PCS_CH0_TX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH0_TX_GEAR_TCLK_SEL                 ("PMA_TCLK"                    ), 
    .PCS_CH0_TX_TCLK2FABRIC_SEL               ("TRUE"                        ), 
    .PCS_CH0_TX_OUTZZ                         ("FALSE"                       ), 
    .PCS_CH0_ENC_DUAL                         ("TRUE"                        ), 
    .PCS_CH0_TX_BITSLIP_DATA_MODE             ("X10"                         ), 
    .PCS_CH0_TX_BRIDGE_CLK_POLINV             ("TX_BRIDGE_CLK"               ),   
    .PCS_CH0_COMMA_REG1                       (10'b1111111111                ), 
    .PCS_CH0_RAPID_IMAX                       (5                             ), 
    .PCS_CH0_RAPID_VMIN_1                     (250                           ), 
    .PCS_CH0_RAPID_VMIN_2                     (1                             ), 
    .PCS_CH0_RX_PRBS_MODE                     ("DISABLE"                     ),            
    .PCS_CH0_RX_ERRCNT_CLR                    ("FALSE"                       ),           
    .PCS_CH0_RX_PRBS_ERR_LPBK                 ("FALSE"                       ), //
    .PCS_CH0_TX_PRBS_MODE                     ("DISABLE"                     ),            
    .PCS_CH0_TX_INSERT_ER                     ("FALSE"                       ),            
    .PCS_CH0_ENABLE_PRBS_GEN                  ("FALSE"                       ),      
    .PCS_CH0_ERR_CNT                          (0                             ),              
    .PCS_CH0_DEFAULT_RADDR                    (6                             ),          
    .PCS_CH0_MASTER_CHECK_OFFSET              (4                             ), 
    .PCS_CH0_DELAY_SET                        (3                             ), 
    .PCS_CH0_SEACH_OFFSET                     ("80BIT"                       ), 
    .PCS_CH0_CEB_RAPIDLS_MMAX                 (5                             ), 
    .PCS_CH0_CTC_AFULL                        (20                            ),            
    .PCS_CH0_CTC_AEMPTY                       (12                            ),           
    .PCS_CH0_CTC_CONTI_SKP_SET                (0                             ),      
    .PCS_CH0_FAR_LOOP                         ("FALSE"                       ),               
    .PCS_CH0_NEAR_LOOP                        ("FALSE"                       ),                
    .PCS_CH0_REG_TX2RX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH0_REG_TX2RX_SLOOP_EN               ("FALSE"                       ), 
    .PCS_CH0_REG_RX2TX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH0_INT_RX_MASK_0                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_1                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_2                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_3                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_4                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_5                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_6                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_MASK_7                    ("FALSE"                       ),          
    .PCS_CH0_INT_RX_CLR_0                     ("FALSE"                       ),             
    .PCS_CH0_INT_RX_CLR_1                     ("FALSE"                       ),             
    .PCS_CH0_INT_RX_CLR_2                     ("FALSE"                       ),             
    .PCS_CH0_INT_RX_CLR_3                     ("FALSE"                       ),             
    .PCS_CH0_INT_RX_CLR_4                     ("FALSE"                       ),           
    .PCS_CH0_INT_RX_CLR_5                     ("FALSE"                       ),           
    .PCS_CH0_INT_RX_CLR_6                     ("FALSE"                       ),           
    .PCS_CH0_INT_RX_CLR_7                     ("FALSE"                       ),            
    .PCS_CH0_CA_RSTN_RX                       ("FALSE"                       ), 
    .PCS_CH0_CA_DYN_DLY_EN_RX                 ("FALSE"                       ), 
    .PCS_CH0_CA_DYN_DLY_SEL_RX                ("FALSE"                       ),
    .PCS_CH0_CA_RX                            (0                             ),
    .PCS_CH0_CA_RSTN_TX                       ("FALSE"                       ), 
    .PCS_CH0_CA_DYN_DLY_EN_TX                 ("FALSE"                       ),    
    .PCS_CH0_CA_DYN_DLY_SEL_TX                ("FALSE"                       ), 
    .PCS_CH0_CA_TX                            (0                             ),    
    .PCS_CH0_RXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_WDALIGN_PWR_REDUCTION            ("NORMAL"                      ), 
    .PCS_CH0_RXDEC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH0_RXCB_PWR_REDUCTION               ("NORMAL"                      ), 
    .PCS_CH0_RXCTC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH0_RXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_RXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH0_RXTEST_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_TXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH0_TXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_TXENC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH0_TXBSLP_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_TXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH0_TXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH0_TXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH0_RXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH0_RXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH0_CTC_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH0_CTC_EMPTY_CHK_EN                 ("TRUE"                        ),
    .PCS_CH0_CEB_FULL_CHK_EN                  ("FALSE"                       ),
    .PCS_CH0_CEB_EMPTY_CHK_EN                 ("FALSE"                       ),
    .PCS_CH0_FLP_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH0_FLP_EMPTY_CHK_EN                 ("TRUE"                        ),  
    .PCS_CH1_BYPASS_WORD_ALIGN                ("TRUE"                        ), 
    .PCS_CH1_BYPASS_DENC                      ("TRUE"                        ), 
    .PCS_CH1_BYPASS_BONDING                   ("TRUE"                        ), 
    .PCS_CH1_BYPASS_CTC                       ("TRUE"                        ), 
    .PCS_CH1_BYPASS_GEAR                      ("FALSE"                       ), 
    .PCS_CH1_BYPASS_BRIDGE                    ("FALSE"                       ), 
    .PCS_CH1_BYPASS_BRIDGE_FIFO               ("FALSE"                       ), 
    .PCS_CH1_DATA_MODE                        ("X16"                         ), 
    .PCS_CH1_RX_POLARITY_INV                  ("DELAY"                       ),            
    .PCS_CH1_ALIGN_MODE                       ("1GB"                         ), 
    .PCS_CH1_SAMP_16B                         ("X16"                         ), 
    .PCS_CH1_FARLP_PWR_REDUCTION              ("FALSE"                       ), 
    .PCS_CH1_COMMA_REG0                       (10'b0000000000                ), 
    .PCS_CH1_COMMA_MASK                       (10'b0                         ), 
    .PCS_CH1_CEB_MODE                         ("10GB"                        ), 
    .PCS_CH1_CTC_MODE                         ("1SKIP"                       ), 
    .PCS_CH1_A_REG                            (8'b01111100                   ), 
    .PCS_CH1_GE_AUTO_EN                       ("FALSE"                       ), 
    .PCS_CH1_SKIP_REG0                        (10'b0                         ), 
    .PCS_CH1_SKIP_REG1                        (10'b0                         ), 
    .PCS_CH1_SKIP_REG2                        (10'b0                         ), 
    .PCS_CH1_SKIP_REG3                        (10'b0                         ), 
    .PCS_CH1_DEC_DUAL                         ("FALSE"                       ), 
    .PCS_CH1_SPLIT                            ("FALSE"                       ), 
    .PCS_CH1_FIFOFLAG_CTC                     ("FALSE"                       ),             
    .PCS_CH1_COMMA_DET_MODE                   ("COMMA_PATTERN"               ), 
    .PCS_CH1_ERRDETECT_SILENCE                ("TRUE"                        ),      
    .PCS_CH1_PMA_RCLK_POLINV                  ("PMA_RCLK"                    ),          
    .PCS_CH1_PCS_RCLK_SEL                     ("PMA_RCLK"                    ), 
    .PCS_CH1_CB_RCLK_SEL                      ("PMA_RCLK"                    ), 
    .PCS_CH1_AFTER_CTC_RCLK_SEL               ("PMA_RCLK"                    ), 
    .PCS_CH1_RCLK_POLINV                      ("RCLK"                        ),            
    .PCS_CH1_BRIDGE_RCLK_SEL                  ("PMA_RCLK"                    ),          
    .PCS_CH1_PCS_RCLK_EN                      ("FALSE"                       ), 
    .PCS_CH1_CB_RCLK_EN                       ("FALSE"                       ), 
    .PCS_CH1_AFTER_CTC_RCLK_EN                ("FALSE"                       ), 
    .PCS_CH1_AFTER_CTC_RCLK_EN_GB             ("TRUE"                        ), 
    .PCS_CH1_AFTER_CTC_RCLK_SEL_1             ("PMA_RCLK"                    ), 
    .PCS_CH1_PCS_RX_RSTN                      ("TRUE"                        ),               
    .PCS_CH1_SLAVE                            ("MASTER"                      ), 
    .PCS_CH1_PCIE_SLAVE                       ("MASTER"                      ), 
    .PCS_CH1_RX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH1_RX_BRIDGE_CLK_POLINV             ("RX_BRIDGE_CLK"               ), 
    .PCS_CH1_AFTER_CTC_RCLK_EN_GB_1           ("TRUE"                        ), 
    .PCS_CH1_PCS_CB_RSTN                      ("TRUE"                        ),               
    .PCS_CH1_TX_BRIDGE_GEAR_SEL               ("FALSE"                       ), 
    .PCS_CH1_TX_BYPASS_BRIDGE_UINT            ("FALSE"                       ), 
    .PCS_CH1_TX_BYPASS_BRIDGE_FIFO            ("FALSE"                       ), 
    .PCS_CH1_TX_BYPASS_GEAR                   ("FALSE"                       ), 
    .PCS_CH1_TX_BYPASS_ENC                    ("TRUE"                        ), 
    .PCS_CH1_TX_BYPASS_BIT_SLIP               ("TRUE"                        ),        
    .PCS_CH1_TX_GEAR_SPLIT                    ("TRUE"                        ), 
    .PCS_CH1_TX_DRIVE_REG_MODE                ("NO_CHANGE"                   ),       
    .PCS_CH1_TX_BIT_SLIP_CYCLES               (0                             ),      
    .PCS_CH1_INT_TX_MASK_0                    ("FALSE"                       ),           
    .PCS_CH1_INT_TX_MASK_1                    ("FALSE"                       ),           
    .PCS_CH1_INT_TX_MASK_2                    ("FALSE"                       ),           
    .PCS_CH1_INT_TX_CLR_0                     ("FALSE"                       ),            
    .PCS_CH1_INT_TX_CLR_1                     ("FALSE"                       ),            
    .PCS_CH1_INT_TX_CLR_2                     ("FALSE"                       ),            
    .PCS_CH1_TX_PMA_TCLK_POLINV               ("PMA_TCLK"                    ),        
    .PCS_CH1_TX_PCS_CLK_EN_SEL                ("TRUE"                        ), 
    .PCS_CH1_TX_BRIDGE_TCLK_SEL               ("TCLK"                        ), 
    .PCS_CH1_TX_TCLK_POLINV                   ("TCLK"                        ),             
    .PCS_CH1_TX_PCS_TCLK_SEL                  ("PMA_TCLK"                    ), 
    .PCS_CH1_TX_PCS_TX_RSTN                   ("TRUE"                        ),             
    .PCS_CH1_TX_SLAVE                         ("MASTER"                      ), 
    .PCS_CH1_TX_GEAR_TCLK_EN_SEL              ("FALSE"                       ), 
    .PCS_CH1_DATA_WIDTH_MODE                  ("X16"                         ), 
    .PCS_CH1_TX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH1_TX_GEAR_TCLK_SEL                 ("PMA_TCLK"                    ), 
    .PCS_CH1_TX_TCLK2FABRIC_SEL               ("TRUE"                        ), 
    .PCS_CH1_TX_OUTZZ                         ("FALSE"                       ), 
    .PCS_CH1_ENC_DUAL                         ("TRUE"                        ), 
    .PCS_CH1_TX_BITSLIP_DATA_MODE             ("X10"                         ),     
    .PCS_CH1_TX_BRIDGE_CLK_POLINV             ("TX_BRIDGE_CLK"               ), 
    .PCS_CH1_COMMA_REG1                       (10'b1111111111                ), 
    .PCS_CH1_RAPID_IMAX                       (5                             ), 
    .PCS_CH1_RAPID_VMIN_1                     (250                           ), 
    .PCS_CH1_RAPID_VMIN_2                     (1                             ), 
    .PCS_CH1_RX_PRBS_MODE                     ("DISABLE"                     ),             
    .PCS_CH1_RX_ERRCNT_CLR                    ("FALSE"                       ),            
    .PCS_CH1_RX_PRBS_ERR_LPBK                 ("FALSE"                       ), 
    .PCS_CH1_TX_PRBS_MODE                     ("DISABLE"                     ),             
    .PCS_CH1_TX_INSERT_ER                     ("FALSE"                       ),             
    .PCS_CH1_ENABLE_PRBS_GEN                  ("FALSE"                       ),          
    .PCS_CH1_ERR_CNT                          (0                             ),                  
    .PCS_CH1_DEFAULT_RADDR                    (6                             ),              
    .PCS_CH1_MASTER_CHECK_OFFSET              (4                             ), 
    .PCS_CH1_DELAY_SET                        (2                             ), 
    .PCS_CH1_SEACH_OFFSET                     ("80BIT"                       ), 
    .PCS_CH1_CEB_RAPIDLS_MMAX                 (5                             ), 
    .PCS_CH1_CTC_AFULL                        (20                            ),                
    .PCS_CH1_CTC_AEMPTY                       (12                            ),               
    .PCS_CH1_CTC_CONTI_SKP_SET                (0                             ),        
    .PCS_CH1_FAR_LOOP                         ("FALSE"                       ),                 
    .PCS_CH1_NEAR_LOOP                        ("FALSE"                       ),                  
    .PCS_CH1_REG_TX2RX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH1_REG_TX2RX_SLOOP_EN               ("FALSE"                       ), 
    .PCS_CH1_REG_RX2TX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH1_INT_RX_MASK_0                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_1                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_2                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_3                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_4                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_5                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_6                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_MASK_7                    ("FALSE"                       ),         
    .PCS_CH1_INT_RX_CLR_0                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_1                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_2                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_3                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_4                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_5                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_6                     ("FALSE"                       ),          
    .PCS_CH1_INT_RX_CLR_7                     ("FALSE"                       ),          
    .PCS_CH1_CA_RSTN_RX                       ("FALSE"                       ), 
    .PCS_CH1_CA_DYN_DLY_EN_RX                 ("FALSE"                       ), 
    .PCS_CH1_CA_DYN_DLY_SEL_RX                ("FALSE"                       ),
    .PCS_CH1_CA_RX                            (0                             ),
    .PCS_CH1_CA_RSTN_TX                       ("FALSE"                       ), 
    .PCS_CH1_CA_DYN_DLY_EN_TX                 ("FALSE"                       ),    
    .PCS_CH1_CA_DYN_DLY_SEL_TX                ("FALSE"                       ), 
    .PCS_CH1_CA_TX                            (0                             ), 
    .PCS_CH1_RXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_WDALIGN_PWR_REDUCTION            ("NORMAL"                      ), 
    .PCS_CH1_RXDEC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH1_RXCB_PWR_REDUCTION               ("NORMAL"                      ), 
    .PCS_CH1_RXCTC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH1_RXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_RXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH1_RXTEST_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_TXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH1_TXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_TXENC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH1_TXBSLP_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_TXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH1_TXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH1_TXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH1_RXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH1_RXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH1_CTC_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH1_CTC_EMPTY_CHK_EN                 ("TRUE"                        ),
    .PCS_CH1_CEB_FULL_CHK_EN                  ("FALSE"                       ),
    .PCS_CH1_CEB_EMPTY_CHK_EN                 ("FALSE"                       ),
    .PCS_CH1_FLP_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH1_FLP_EMPTY_CHK_EN                 ("TRUE"                        ),  
    .PCS_CH2_BYPASS_WORD_ALIGN                ("FALSE"                       ), 
    .PCS_CH2_BYPASS_DENC                      ("FALSE"                       ), 
    .PCS_CH2_BYPASS_BONDING                   ("TRUE"                        ), 
    .PCS_CH2_BYPASS_CTC                       ("TRUE"                        ), 
    .PCS_CH2_BYPASS_GEAR                      ("FALSE"                       ), 
    .PCS_CH2_BYPASS_BRIDGE                    ("FALSE"                       ), 
    .PCS_CH2_BYPASS_BRIDGE_FIFO               ("FALSE"                       ), 
    .PCS_CH2_DATA_MODE                        ("X20"                         ), 
    .PCS_CH2_RX_POLARITY_INV                  ("DELAY"                       ),        
    .PCS_CH2_ALIGN_MODE                       ("1GB"                         ), 
    .PCS_CH2_SAMP_16B                         ("X20"                         ), 
    .PCS_CH2_FARLP_PWR_REDUCTION              ("FALSE"                       ), 
    .PCS_CH2_COMMA_REG0                       (10'b0101111100                ), 
    .PCS_CH2_COMMA_MASK                       (10'b0000000000                ), 
    .PCS_CH2_CEB_MODE                         ("10GB"                        ), 
    .PCS_CH2_CTC_MODE                         ("1SKIP"                       ), 
    .PCS_CH2_A_REG                            (8'b01111100                   ), 
    .PCS_CH2_GE_AUTO_EN                       ("FALSE"                       ), 
    .PCS_CH2_SKIP_REG0                        (10'b0                         ), 
    .PCS_CH2_SKIP_REG1                        (10'b0                         ), 
    .PCS_CH2_SKIP_REG2                        (10'b0                         ), 
    .PCS_CH2_SKIP_REG3                        (10'b0                         ), 
    .PCS_CH2_DEC_DUAL                         ("TRUE"                        ), 
    .PCS_CH2_SPLIT                            ("FALSE"                       ), 
    .PCS_CH2_FIFOFLAG_CTC                     ("FALSE"                       ),           
    .PCS_CH2_COMMA_DET_MODE                   ("COMMA_PATTERN"               ), 
    .PCS_CH2_ERRDETECT_SILENCE                ("TRUE"                        ),    
    .PCS_CH2_PMA_RCLK_POLINV                  ("PMA_RCLK"                    ),        
    .PCS_CH2_PCS_RCLK_SEL                     ("PMA_RCLK"                    ), 
    .PCS_CH2_CB_RCLK_SEL                      ("PMA_RCLK"                    ), 
    .PCS_CH2_AFTER_CTC_RCLK_SEL               ("PMA_RCLK"                    ), 
    .PCS_CH2_RCLK_POLINV                      ("RCLK"                        ),          
    .PCS_CH2_BRIDGE_RCLK_SEL                  ("PMA_RCLK"                    ),        
    .PCS_CH2_PCS_RCLK_EN                      ("FALSE"                       ), 
    .PCS_CH2_CB_RCLK_EN                       ("FALSE"                       ), 
    .PCS_CH2_AFTER_CTC_RCLK_EN                ("FALSE"                       ), 
    .PCS_CH2_AFTER_CTC_RCLK_EN_GB             ("TRUE"                        ), 
    .PCS_CH2_AFTER_CTC_RCLK_SEL_1             ("PMA_RCLK"                    ), 
    .PCS_CH2_PCS_RX_RSTN                      ("TRUE"                        ),            
    .PCS_CH2_SLAVE                            ("MASTER"                      ), 
    .PCS_CH2_PCIE_SLAVE                       ("MASTER"                      ), 
    .PCS_CH2_RX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH2_RX_BRIDGE_CLK_POLINV             ("RX_BRIDGE_CLK"               ), 
    .PCS_CH2_AFTER_CTC_RCLK_EN_GB_1           ("TRUE"                        ), 
    .PCS_CH2_PCS_CB_RSTN                      ("TRUE"                        ),            
    .PCS_CH2_TX_BRIDGE_GEAR_SEL               ("FALSE"                       ), 
    .PCS_CH2_TX_BYPASS_BRIDGE_UINT            ("FALSE"                       ), 
    .PCS_CH2_TX_BYPASS_BRIDGE_FIFO            ("FALSE"                       ), 
    .PCS_CH2_TX_BYPASS_GEAR                   ("FALSE"                       ), 
    .PCS_CH2_TX_BYPASS_ENC                    ("FALSE"                       ), 
    .PCS_CH2_TX_BYPASS_BIT_SLIP               ("TRUE"                        ),     
    .PCS_CH2_TX_GEAR_SPLIT                    ("TRUE"                        ), 
    .PCS_CH2_TX_DRIVE_REG_MODE                ("NO_CHANGE"                   ),    
    .PCS_CH2_TX_BIT_SLIP_CYCLES               (0                             ),   
    .PCS_CH2_INT_TX_MASK_0                    ("FALSE"                       ),        
    .PCS_CH2_INT_TX_MASK_1                    ("FALSE"                       ),        
    .PCS_CH2_INT_TX_MASK_2                    ("FALSE"                       ),          
    .PCS_CH2_INT_TX_CLR_0                     ("FALSE"                       ),           
    .PCS_CH2_INT_TX_CLR_1                     ("FALSE"                       ),           
    .PCS_CH2_INT_TX_CLR_2                     ("FALSE"                       ),                
    .PCS_CH2_TX_PMA_TCLK_POLINV               ("PMA_TCLK"                    ),       
    .PCS_CH2_TX_PCS_CLK_EN_SEL                ("TRUE"                        ), 
    .PCS_CH2_TX_BRIDGE_TCLK_SEL               ("TCLK"                        ), 
    .PCS_CH2_TX_TCLK_POLINV                   ("TCLK"                        ),             
    .PCS_CH2_TX_PCS_TCLK_SEL                  ("PMA_TCLK"                    ), 
    .PCS_CH2_TX_PCS_TX_RSTN                   ("TRUE"                        ),           
    .PCS_CH2_TX_SLAVE                         ("MASTER"                      ), 
    .PCS_CH2_TX_GEAR_TCLK_EN_SEL              ("FALSE"                       ), 
    .PCS_CH2_DATA_WIDTH_MODE                  ("X20"                         ), 
    .PCS_CH2_TX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH2_TX_GEAR_TCLK_SEL                 ("PMA_TCLK"                    ), 
    .PCS_CH2_TX_TCLK2FABRIC_SEL               ("TRUE"                        ), 
    .PCS_CH2_TX_OUTZZ                         ("FALSE"                       ), 
    .PCS_CH2_ENC_DUAL                         ("TRUE"                        ), 
    .PCS_CH2_TX_BITSLIP_DATA_MODE             ("X10"                         ),      
    .PCS_CH2_TX_BRIDGE_CLK_POLINV             ("TX_BRIDGE_CLK"               ), 
    .PCS_CH2_COMMA_REG1                       (10'b1010000011                ), 
    .PCS_CH2_RAPID_IMAX                       (5                             ), 
    .PCS_CH2_RAPID_VMIN_1                     (250                           ), 
    .PCS_CH2_RAPID_VMIN_2                     (1                             ), 
    .PCS_CH2_RX_PRBS_MODE                     ("DISABLE"                     ),            
    .PCS_CH2_RX_ERRCNT_CLR                    ("FALSE"                       ),           
    .PCS_CH2_RX_PRBS_ERR_LPBK                 ("FALSE"                       ), 
    .PCS_CH2_TX_PRBS_MODE                     ("DISABLE"                     ),             
    .PCS_CH2_TX_INSERT_ER                     ("FALSE"                       ),            
    .PCS_CH2_ENABLE_PRBS_GEN                  ("FALSE"                       ),          
    .PCS_CH2_ERR_CNT                          (0                             ),                 
    .PCS_CH2_DEFAULT_RADDR                    (6                             ),              
    .PCS_CH2_MASTER_CHECK_OFFSET              (4                             ), 
    .PCS_CH2_DELAY_SET                        (1                             ), 
    .PCS_CH2_SEACH_OFFSET                     ("80BIT"                       ), 
    .PCS_CH2_CEB_RAPIDLS_MMAX                 (5                             ), 
    .PCS_CH2_CTC_AFULL                        (20                            ),            
    .PCS_CH2_CTC_AEMPTY                       (12                            ),            
    .PCS_CH2_CTC_CONTI_SKP_SET                (0                             ),      
    .PCS_CH2_FAR_LOOP                         ("FALSE"                       ),                        
    .PCS_CH2_NEAR_LOOP                        ("FALSE"                       ),                
    .PCS_CH2_REG_TX2RX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH2_REG_TX2RX_SLOOP_EN               ("FALSE"                       ), 
    .PCS_CH2_REG_RX2TX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH2_INT_RX_MASK_0                    ("FALSE"                       ),         
    .PCS_CH2_INT_RX_MASK_1                    ("FALSE"                       ),          
    .PCS_CH2_INT_RX_MASK_2                    ("FALSE"                       ),         
    .PCS_CH2_INT_RX_MASK_3                    ("FALSE"                       ),        
    .PCS_CH2_INT_RX_MASK_4                    ("FALSE"                       ),             
    .PCS_CH2_INT_RX_MASK_5                    ("FALSE"                       ),             
    .PCS_CH2_INT_RX_MASK_6                    ("FALSE"                       ),             
    .PCS_CH2_INT_RX_MASK_7                    ("FALSE"                       ),                 
    .PCS_CH2_INT_RX_CLR_0                     ("FALSE"                       ),           
    .PCS_CH2_INT_RX_CLR_1                     ("FALSE"                       ),               
    .PCS_CH2_INT_RX_CLR_2                     ("FALSE"                       ),          
    .PCS_CH2_INT_RX_CLR_3                     ("FALSE"                       ),         
    .PCS_CH2_INT_RX_CLR_4                     ("FALSE"                       ),         
    .PCS_CH2_INT_RX_CLR_5                     ("FALSE"                       ),             
    .PCS_CH2_INT_RX_CLR_6                     ("FALSE"                       ),             
    .PCS_CH2_INT_RX_CLR_7                     ("FALSE"                       ),            
    .PCS_CH2_CA_RSTN_RX                       ("FALSE"                       ), 
    .PCS_CH2_CA_DYN_DLY_EN_RX                 ("FALSE"                       ), 
    .PCS_CH2_CA_DYN_DLY_SEL_RX                ("FALSE"                       ),
    .PCS_CH2_CA_RX                            (0                             ),
    .PCS_CH2_CA_RSTN_TX                       ("FALSE"                       ), 
    .PCS_CH2_CA_DYN_DLY_EN_TX                 ("FALSE"                       ),    
    .PCS_CH2_CA_DYN_DLY_SEL_TX                ("FALSE"                       ), 
    .PCS_CH2_CA_TX                            (0                             ), 
    .PCS_CH2_RXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_WDALIGN_PWR_REDUCTION            ("NORMAL"                      ), 
    .PCS_CH2_RXDEC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH2_RXCB_PWR_REDUCTION               ("NORMAL"                      ), 
    .PCS_CH2_RXCTC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH2_RXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_RXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH2_RXTEST_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_TXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH2_TXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_TXENC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH2_TXBSLP_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_TXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH2_TXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH2_TXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH2_RXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH2_RXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH2_CTC_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH2_CTC_EMPTY_CHK_EN                 ("TRUE"                        ),
    .PCS_CH2_CEB_FULL_CHK_EN                  ("FALSE"                       ),
    .PCS_CH2_CEB_EMPTY_CHK_EN                 ("FALSE"                       ),
    .PCS_CH2_FLP_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH2_FLP_EMPTY_CHK_EN                 ("TRUE"                        ),  
    .PCS_CH3_BYPASS_WORD_ALIGN                ("FALSE"                       ), 
    .PCS_CH3_BYPASS_DENC                      ("FALSE"                       ), 
    .PCS_CH3_BYPASS_BONDING                   ("TRUE"                        ), 
    .PCS_CH3_BYPASS_CTC                       ("TRUE"                        ), 
    .PCS_CH3_BYPASS_GEAR                      ("FALSE"                       ), 
    .PCS_CH3_BYPASS_BRIDGE                    ("FALSE"                       ), 
    .PCS_CH3_BYPASS_BRIDGE_FIFO               ("FALSE"                       ), 
    .PCS_CH3_DATA_MODE                        ("X20"                         ), 
    .PCS_CH3_RX_POLARITY_INV                  ("DELAY"                       ),         
    .PCS_CH3_ALIGN_MODE                       ("10GB"                        ), 
    .PCS_CH3_SAMP_16B                         ("X20"                         ), 
    .PCS_CH3_FARLP_PWR_REDUCTION              ("FALSE"                       ), 
    .PCS_CH3_COMMA_REG0                       (10'b0101111100                ), 
    .PCS_CH3_COMMA_MASK                       (10'b1110000000                ), 
    .PCS_CH3_CEB_MODE                         ("10GB"                        ), 
    .PCS_CH3_CTC_MODE                         ("1SKIP"                       ), 
    .PCS_CH3_A_REG                            (8'b01111100                   ), 
    .PCS_CH3_GE_AUTO_EN                       ("FALSE"                       ), 
    .PCS_CH3_SKIP_REG0                        (10'b0                         ), 
    .PCS_CH3_SKIP_REG1                        (10'b0                         ), 
    .PCS_CH3_SKIP_REG2                        (10'b0                         ), 
    .PCS_CH3_SKIP_REG3                        (10'b0                         ), 
    .PCS_CH3_DEC_DUAL                         ("TRUE"                        ), 
    .PCS_CH3_SPLIT                            ("FALSE"                       ), 
    .PCS_CH3_FIFOFLAG_CTC                     ("FALSE"                       ),           
    .PCS_CH3_COMMA_DET_MODE                   ("COMMA_PATTERN"               ), 
    .PCS_CH3_ERRDETECT_SILENCE                ("TRUE"                        ),       
    .PCS_CH3_PMA_RCLK_POLINV                  ("PMA_RCLK"                    ),            
    .PCS_CH3_PCS_RCLK_SEL                     ("PMA_RCLK"                    ), 
    .PCS_CH3_CB_RCLK_SEL                      ("PMA_RCLK"                    ), 
    .PCS_CH3_AFTER_CTC_RCLK_SEL               ("PMA_RCLK"                    ), 
    .PCS_CH3_RCLK_POLINV                      ("RCLK"                        ),           
    .PCS_CH3_BRIDGE_RCLK_SEL                  ("PMA_RCLK"                    ),         
    .PCS_CH3_PCS_RCLK_EN                      ("FALSE"                       ), 
    .PCS_CH3_CB_RCLK_EN                       ("FALSE"                       ), 
    .PCS_CH3_AFTER_CTC_RCLK_EN                ("FALSE"                       ), 
    .PCS_CH3_AFTER_CTC_RCLK_EN_GB             ("TRUE"                        ), 
    .PCS_CH3_AFTER_CTC_RCLK_SEL_1             ("PMA_RCLK"                    ), 
    .PCS_CH3_PCS_RX_RSTN                      ("TRUE"                        ),               
    .PCS_CH3_SLAVE                            ("MASTER"                      ), 
    .PCS_CH3_PCIE_SLAVE                       ("MASTER"                      ), 
    .PCS_CH3_RX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH3_RX_BRIDGE_CLK_POLINV             ("RX_BRIDGE_CLK"               ), 
    .PCS_CH3_AFTER_CTC_RCLK_EN_GB_1           ("TRUE"                        ), 
    .PCS_CH3_PCS_CB_RSTN                      ("TRUE"                        ),             
    .PCS_CH3_TX_BRIDGE_GEAR_SEL               ("FALSE"                       ), 
    .PCS_CH3_TX_BYPASS_BRIDGE_UINT            ("FALSE"                       ), 
    .PCS_CH3_TX_BYPASS_BRIDGE_FIFO            ("FALSE"                       ), 
    .PCS_CH3_TX_BYPASS_GEAR                   ("FALSE"                       ), 
    .PCS_CH3_TX_BYPASS_ENC                    ("FALSE"                       ), 
    .PCS_CH3_TX_BYPASS_BIT_SLIP               ("TRUE"                        ),         
    .PCS_CH3_TX_GEAR_SPLIT                    ("TRUE"                        ), 
    .PCS_CH3_TX_DRIVE_REG_MODE                ("NO_CHANGE"                   ),         
    .PCS_CH3_TX_BIT_SLIP_CYCLES               (0                             ),      
    .PCS_CH3_INT_TX_MASK_0                    ("FALSE"                       ),        
    .PCS_CH3_INT_TX_MASK_1                    ("FALSE"                       ),        
    .PCS_CH3_INT_TX_MASK_2                    ("FALSE"                       ),        
    .PCS_CH3_INT_TX_CLR_0                     ("FALSE"                       ),         
    .PCS_CH3_INT_TX_CLR_1                     ("FALSE"                       ),         
    .PCS_CH3_INT_TX_CLR_2                     ("FALSE"                       ),         
    .PCS_CH3_TX_PMA_TCLK_POLINV               ("PMA_TCLK"                    ),          
    .PCS_CH3_TX_PCS_CLK_EN_SEL                ("TRUE"                        ), 
    .PCS_CH3_TX_BRIDGE_TCLK_SEL               ("TCLK"                        ), 
    .PCS_CH3_TX_TCLK_POLINV                   ("TCLK"                        ),              
    .PCS_CH3_TX_PCS_TCLK_SEL                  ("PMA_TCLK"                    ), 
    .PCS_CH3_TX_PCS_TX_RSTN                   ("TRUE"                        ),              
    .PCS_CH3_TX_SLAVE                         ("MASTER"                      ), 
    .PCS_CH3_TX_GEAR_TCLK_EN_SEL              ("FALSE"                       ), 
    .PCS_CH3_DATA_WIDTH_MODE                  ("X20"                         ), 
    .PCS_CH3_TX_64B66B_67B                    ("NORMAL"                      ), 
    .PCS_CH3_TX_GEAR_TCLK_SEL                 ("PMA_TCLK"                    ), 
    .PCS_CH3_TX_TCLK2FABRIC_SEL               ("TRUE"                        ), 
    .PCS_CH3_TX_OUTZZ                         ("FALSE"                       ), 
    .PCS_CH3_ENC_DUAL                         ("TRUE"                        ), 
    .PCS_CH3_TX_BITSLIP_DATA_MODE             ("X10"                         ),      
    .PCS_CH3_TX_BRIDGE_CLK_POLINV             ("TX_BRIDGE_CLK"               ), 
    .PCS_CH3_COMMA_REG1                       (10'b1010000011                ), 
    .PCS_CH3_RAPID_IMAX                       (5                             ), 
    .PCS_CH3_RAPID_VMIN_1                     (250                           ), 
    .PCS_CH3_RAPID_VMIN_2                     (1                             ), 
    .PCS_CH3_RX_PRBS_MODE                     ("DISABLE"                     ),             
    .PCS_CH3_RX_ERRCNT_CLR                    ("FALSE"                       ),            
    .PCS_CH3_RX_PRBS_ERR_LPBK                 ("FALSE"                       ), 
    .PCS_CH3_TX_PRBS_MODE                     ("DISABLE"                     ),             
    .PCS_CH3_TX_INSERT_ER                     ("FALSE"                       ),             
    .PCS_CH3_ENABLE_PRBS_GEN                  ("FALSE"                       ),          
    .PCS_CH3_ERR_CNT                          (0                             ),                  
    .PCS_CH3_DEFAULT_RADDR                    (6                             ),               
    .PCS_CH3_MASTER_CHECK_OFFSET              (4                             ), 
    .PCS_CH3_DELAY_SET                        (0                             ), 
    .PCS_CH3_SEACH_OFFSET                     ("80BIT"                       ), 
    .PCS_CH3_CEB_RAPIDLS_MMAX                 (5                             ), 
    .PCS_CH3_CTC_AFULL                        (20                            ),                 
    .PCS_CH3_CTC_AEMPTY                       (12                            ),                
    .PCS_CH3_CTC_CONTI_SKP_SET                (0                             ),         
    .PCS_CH3_FAR_LOOP                         ("FALSE"                       ),                  
    .PCS_CH3_NEAR_LOOP                        ("FALSE"                       ),                   
    .PCS_CH3_REG_TX2RX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH3_REG_TX2RX_SLOOP_EN               ("FALSE"                       ), 
    .PCS_CH3_REG_RX2TX_PLOOP_EN               ("FALSE"                       ), 
    .PCS_CH3_INT_RX_MASK_0                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_1                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_2                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_3                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_4                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_5                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_6                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_MASK_7                    ("FALSE"                       ),             
    .PCS_CH3_INT_RX_CLR_0                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_1                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_2                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_3                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_4                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_5                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_6                     ("FALSE"                       ),              
    .PCS_CH3_INT_RX_CLR_7                     ("FALSE"                       ),              
    .PCS_CH3_CA_RSTN_RX                       ("FALSE"                       ), 
    .PCS_CH3_CA_DYN_DLY_EN_RX                 ("FALSE"                       ), 
    .PCS_CH3_CA_DYN_DLY_SEL_RX                ("FALSE"                       ),
    .PCS_CH3_CA_RX                            (0                             ),
    .PCS_CH3_CA_RSTN_TX                       ("FALSE"                       ), 
    .PCS_CH3_CA_DYN_DLY_EN_TX                 ("FALSE"                       ),    
    .PCS_CH3_CA_DYN_DLY_SEL_TX                ("FALSE"                       ), 
    .PCS_CH3_CA_TX                            (0                             ), 
    .PCS_CH3_RXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_WDALIGN_PWR_REDUCTION            ("NORMAL"                      ), 
    .PCS_CH3_RXDEC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH3_RXCB_PWR_REDUCTION               ("NORMAL"                      ), 
    .PCS_CH3_RXCTC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH3_RXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_RXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH3_RXTEST_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_TXBRG_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH3_TXGEAR_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_TXENC_PWR_REDUCTION              ("NORMAL"                      ), 
    .PCS_CH3_TXBSLP_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_TXPRBS_PWR_REDUCTION             ("NORMAL"                      ), 
    .PCS_CH3_TXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH3_TXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH3_RXBRG_FULL_CHK_EN                ("FALSE"                       ),
    .PCS_CH3_RXBRG_EMPTY_CHK_EN               ("FALSE"                       ),
    .PCS_CH3_CTC_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH3_CTC_EMPTY_CHK_EN                 ("TRUE"                        ),
    .PCS_CH3_CEB_FULL_CHK_EN                  ("FALSE"                       ),
    .PCS_CH3_CEB_EMPTY_CHK_EN                 ("FALSE"                       ),
    .PCS_CH3_FLP_FULL_CHK_EN                  ("TRUE"                        ),
    .PCS_CH3_FLP_EMPTY_CHK_EN                 ("TRUE"                        ),
    .PMA_CH0_REG_RX_PD                        ("ON"                          ),                  
    .PMA_CH0_REG_RX_PD_EN                     ("FALSE"                       ),              
    .PMA_CH0_REG_RX_CLKPATH_PD                ("ON"                          ),         
    .PMA_CH0_REG_RX_CLKPATH_PD_EN             ("FALSE"                       ),      
    .PMA_CH0_REG_RX_DATAPATH_PD               ("ON"                          ),        
    .PMA_CH0_REG_RX_DATAPATH_PD_EN            ("FALSE"                       ),     
    .PMA_CH0_REG_RX_SIGDET_PD                 ("ON"                          ),          
    .PMA_CH0_REG_RX_SIGDET_PD_EN              ("FALSE"                       ),       
    .PMA_CH0_REG_RX_DCC_RST_N                 ("TRUE"                        ),          
    .PMA_CH0_REG_RX_DCC_RST_N_EN              ("TRUE"                        ),       
    .PMA_CH0_REG_RX_CDR_RST_N                 ("TRUE"                        ),          
    .PMA_CH0_REG_RX_CDR_RST_N_EN              ("FALSE"                       ),       
    .PMA_CH0_REG_RX_SIGDET_RST_N              ("TRUE"                        ),       
    .PMA_CH0_REG_RX_SIGDET_RST_N_EN           ("FALSE"                       ),    
    .PMA_CH0_REG_RXPCLK_SLIP                  ("FALSE"                       ),           
    .PMA_CH0_REG_RXPCLK_SLIP_OW               ("DISABLE"                     ),        
    .PMA_CH0_REG_RX_PCLKSWITCH_RST_N          ("TRUE"                        ),   
    .PMA_CH0_REG_RX_PCLKSWITCH_RST_N_EN       ("FALSE"                       ),
    .PMA_CH0_REG_RX_PCLKSWITCH                ("FALSE"                       ),          
    .PMA_CH0_REG_RX_PCLKSWITCH_EN             ("FALSE"                       ),         
    .PMA_CH0_REG_RX_HIGHZ                     ("FALSE"                       ), 
    .PMA_CH0_REG_RX_HIGHZ_EN                  ("FALSE"                       ), 
    .PMA_CH0_REG_RX_EQ_C_SET                  (0                             ),            
    .PMA_CH0_REG_RX_EQ_R_SET                  (1                             ),              
    .PMA_CH0_REG_RX_BUSWIDTH                  ("16BIT"                       ), 
    .PMA_CH0_REG_RX_BUSWIDTH_EN               ("TRUE"                        ), 
    .PMA_CH0_REG_RX_RATE                      ("DIV4"                        ),                
    .PMA_CH0_REG_RX_RATE_EN                   ("FALSE"                       ),             
    .PMA_CH0_REG_RX_RES_TRIM                  (51                            ),            
    .PMA_CH0_REG_RX_RES_TRIM_EN               ("FALSE"                       ),         
    .PMA_CH0_REG_RX_EQ_OFF                    ("FALSE"                       ),              
    .PMA_CH0_REG_RX_PREAMP_IC                 (1367                          ),           
    .PMA_CH0_REG_RX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),       
    .PMA_CH0_REG_RX_PIBUF_IC                  (2                             ),            
    .PMA_CH0_REG_RX_DCC_IC_RX                 (3                             ),           
    .PMA_CH0_REG_RX_DCC_IC_TX                 (3                             ),           
    .PMA_CH0_REG_RX_ICTRL_TRX                 ("100PCT"                      ),           
    .PMA_CH0_REG_RX_ICTRL_PREAMP              ("100PCT"                      ),        
    .PMA_CH0_REG_RX_ICTRL_SLICER              ("100PCT"                      ),        
    .PMA_CH0_REG_RX_ICTRL_PIBUF               ("100PCT"                      ),         
    .PMA_CH0_REG_RX_ICTRL_PI                  ("100PCT"                      ),            
    .PMA_CH0_REG_RX_ICTRL_DCC                 ("100PCT"                      ),           
    .PMA_CH0_REG_RX_ICTRL_PREDRV              ("100PCT"                      ),         
    .PMA_CH0_REG_TX_RATE                      ("DIV4"                        ),                
    .PMA_CH0_REG_TX_RATE_EN                   ("FALSE"                       ),             
    .PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N         ("TRUE"                        ),   
    .PMA_CH0_REG_RX_TX2RX_PLPBK_RST_N_EN      ("FALSE"                       ),
    .PMA_CH0_REG_RX_TX2RX_PLPBK_EN            ("FALSE"                       ),          
    .PMA_CH0_REG_TXCLK_SEL                    ("PLL"                         ),                  
    .PMA_CH0_REG_RX_DATA_POLARITY             ("NORMAL"                      ),           
    .PMA_CH0_REG_RX_ERR_INSERT                ("FALSE"                       ),             
    .PMA_CH0_REG_UDP_CHK_EN                   ("FALSE"                       ),                 
    .PMA_CH0_REG_PRBS_SEL                     ("PRBS7"                       ),                   
    .PMA_CH0_REG_PRBS_CHK_EN                  ("FALSE"                       ),                 
    .PMA_CH0_REG_PRBS_CHK_WIDTH_SEL           ("16BIT"                       ),           
    .PMA_CH0_REG_BIST_CHK_PAT_SEL             ("PRBS"                        ),           
    .PMA_CH0_REG_LOAD_ERR_CNT                 ("DISABLE"                     ),               
    .PMA_CH0_REG_CHK_COUNTER_EN               ("FALSE"                       ),             
    .PMA_CH0_REG_CDR_PROP_TURBO_GAIN          (6                             ),        
    .PMA_CH0_REG_CDR_INT_GAIN                 (5                             ),               
    .PMA_CH0_REG_CDR_INT_TURBO_GAIN           (6                             ),         
    .PMA_CH0_REG_CDR_INT_SAT_MAX              (992                           ),            
    .PMA_CH0_REG_CDR_INT_SAT_MIN              (32                            ),            
    .PMA_CH0_REG_CDR_INT_RST                  ("FALSE"                       ),                
    .PMA_CH0_REG_CDR_INT_RST_OW               ("DISABLE"                     ),             
    .PMA_CH0_REG_CDR_PROP_RST                 ("FALSE"                       ),               
    .PMA_CH0_REG_CDR_PROP_RST_OW              ("DISABLE"                     ),            
    .PMA_CH0_REG_CDR_LOCK_RST                 ("FALSE"                       ),               
    .PMA_CH0_REG_CDR_LOCK_RST_OW              ("DISABLE"                     ),            
    .PMA_CH0_REG_CDR_RX_PI_FORCE_SEL          (0                             ),        
    .PMA_CH0_REG_CDR_RX_PI_FORCE_D            (0                             ),            
    .PMA_CH0_REG_CDR_LOCK_TIMER               ("25_6U"                       ), 
    .PMA_CH0_REG_CDR_TURBO_MODE_TIMER         (1                             ),       
    .PMA_CH0_REG_CDR_LOCK_VAL                 ("FALSE"                       ),               
    .PMA_CH0_REG_CDR_LOCK_OW                  ("DISABLE"                     ),                
    .PMA_CH0_REG_CDR_INT_SAT_DET_EN           ("TRUE"                        ),         
    .PMA_CH0_REG_CDR_SAT_DET_STATUS_EN        ("FALSE"                       ),      
    .PMA_CH0_REG_CDR_SAT_DET_STATUS_RESET_EN  ("FALSE"                       ),
    .PMA_CH0_REG_CDR_PI_CTRL_RST              ("FALSE"                       ),              
    .PMA_CH0_REG_CDR_PI_CTRL_RST_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_CDR_SAT_DET_RST              ("FALSE"                       ),              
    .PMA_CH0_REG_CDR_SAT_DET_RST_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_CDR_SAT_DET_STICKY_RST       ("FALSE"                       ),       
    .PMA_CH0_REG_CDR_SAT_DET_STICKY_RST_OW    ("DISABLE"                     ),    
    .PMA_CH0_REG_CDR_SIGDET_STATUS_DIS        ("FALSE"                       ),        
    .PMA_CH0_REG_CDR_SAT_DET_TIMER            (2                             ),            
    .PMA_CH0_REG_CDR_SAT_DET_STATUS_VAL       ("FALSE"                       ),       
    .PMA_CH0_REG_CDR_SAT_DET_STATUS_OW        ("DISABLE"                     ),        
    .PMA_CH0_REG_CDR_TURBO_MODE_EN            ("TRUE"                        ),            
    .PMA_CH0_REG_CDR_STATUS_RADDR_INIT        (0                             ),        
    .PMA_CH0_REG_CDR_STATUS_FIFO_EN           ("TRUE"                        ),           
    .PMA_CH0_REG_PMA_TEST_SEL                 (0                             ),                 
    .PMA_CH0_REG_OOB_COMWAKE_GAP_MIN          (3                             ),          
    .PMA_CH0_REG_OOB_COMWAKE_GAP_MAX          (11                            ),          
    .PMA_CH0_REG_OOB_COMINIT_GAP_MIN          (15                            ),          
    .PMA_CH0_REG_OOB_COMINIT_GAP_MAX          (35                            ),          
    .PMA_CH0_REG_RX_PIBUF_IC_TX               (1                             ),               
    .PMA_CH0_REG_COMWAKE_STATUS_CLEAR         (0                             ),         
    .PMA_CH0_REG_COMINIT_STATUS_CLEAR         (0                             ),         
    .PMA_CH0_REG_RX_SYNC_RST_N_EN             ("FALSE"                       ),             
    .PMA_CH0_REG_RX_SYNC_RST_N                ("TRUE"                        ),                
    .PMA_CH0_REG_RX_SATA_COMINIT_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_RX_SATA_COMINIT              ("FALSE"                       ),              
    .PMA_CH0_REG_RX_SATA_COMWAKE_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_RX_SATA_COMWAKE              ("FALSE"                       ),              
    .PMA_CH0_REG_RX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH0_REG_TX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH0_REG_RX_SLIP_SEL_EN               ("FALSE"                       ),               
    .PMA_CH0_REG_RX_SLIP_SEL                  (0                             ),                  
    .PMA_CH0_REG_RX_SLIP_EN                   ("FALSE"                       ),                   
    .PMA_CH0_REG_RX_SIGDET_STATUS_SEL         (5                             ),         
    .PMA_CH0_REG_RX_SIGDET_FSM_RST_N          ("TRUE"                        ),          
    .PMA_CH0_REG_RX_SIGDET_STATUS_OW          ("DISABLE"                     ),          
    .PMA_CH0_REG_RX_SIGDET_STATUS             ("FALSE"                       ),             
    .PMA_CH0_REG_RX_SIGDET_GRM                (0                             ),                
    .PMA_CH0_REG_RX_SIGDET_PULSE_EXT          ("DISABLE"                     ),          
    .PMA_CH0_REG_RX_SIGDET_CH2_SEL            (0                             ),            
    .PMA_CH0_REG_RX_SIGDET_CH2_CHK_WINDOW     (3                             ),     
    .PMA_CH0_REG_RX_SIGDET_CHK_WINDOW_EN      ("TRUE"                        ),      
    .PMA_CH0_REG_RX_SIGDET_NOSIG_COUNT_SETTING(4                             ),
    .PMA_CH0_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (0                             ),  
    .PMA_CH0_REG_SLIP_FIFO_INV_EN             ("FALSE"                       ),             
    .PMA_CH0_REG_SLIP_FIFO_INV                ("POS_EDGE"                    ),                
    .PMA_CH0_REG_RX_SIGDET_4OOB_DET_SEL       (7                             ),       
    .PMA_CH0_REG_RX_SIGDET_IC_I               (10                            ),               
    .PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N_OW   ("DISABLE"                     ),   
    .PMA_CH0_REG_RX_OOB_DETECTOR_RESET_N      ("FALSE"                       ),      
    .PMA_CH0_REG_RX_OOB_DETECTOR_PD_OW        ("DISABLE"                     ),        
    .PMA_CH0_REG_RX_OOB_DETECTOR_PD           ("ON"                          ),           
    .PMA_CH0_REG_RX_TERM_CM_CTRL              ("5DIV7"                       ),              
    .PMA_CH0_REG_TX_PD                        ("ON"                          ),                        
    .PMA_CH0_REG_TX_PD_OW                     ("DISABLE"                     ),                     
    .PMA_CH0_REG_TX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH0_REG_TX_CLKPATH_PD_OW             ("DISABLE"                     ),             
    .PMA_CH0_REG_TX_BEACON_TIMER_SEL          (0                             ),          
    .PMA_CH0_REG_TX_RXDET_REQ_OW              ("DISABLE"                     ),              
    .PMA_CH0_REG_TX_RXDET_REQ                 ("FALSE"                       ),                 
    .PMA_CH0_REG_TX_BEACON_EN_OW              ("DISABLE"                     ),              
    .PMA_CH0_REG_TX_BEACON_EN                 ("FALSE"                       ),                 
    .PMA_CH0_REG_TX_EI_EN_OW                  ("DISABLE"                     ),                  
    .PMA_CH0_REG_TX_EI_EN                     ("FALSE"                       ),                     
    .PMA_CH0_REG_TX_RES_CAL_EN                ("FALSE"                       ),                
    .PMA_CH0_REG_TX_RES_CAL                   (51                            ),                   
    .PMA_CH0_REG_TX_BIAS_CAL_EN               ("FALSE"                       ),               
    .PMA_CH0_REG_TX_BIAS_CTRL                 (48                            ),                 
    .PMA_CH0_REG_TX_RXDET_TIMER_SEL           ("12CYCLE"                     ),           
    .PMA_CH0_REG_TX_SYNC_OW                   ("DISABLE"                     ),                   
    .PMA_CH0_REG_TX_SYNC                      ("DISABLE"                     ),                        
    .PMA_CH0_REG_TX_PD_POST                   ("OFF"                         ), 
    .PMA_CH0_REG_TX_PD_POST_OW                ("ENABLE"                      ),                
    .PMA_CH0_REG_TX_RESET_N_OW                ("DISABLE"                     ),                
    .PMA_CH0_REG_TX_RESET_N                   ("TRUE"                        ),                   
    .PMA_CH0_REG_TX_DCC_RESET_N_OW            ("DISABLE"                     ),            
    .PMA_CH0_REG_TX_DCC_RESET_N               ("TRUE"                        ),                 
    .PMA_CH0_REG_TX_BUSWIDTH_OW               ("ENABLE"                      ), 
    .PMA_CH0_REG_TX_BUSWIDTH                  ("16BIT"                       ), 
    .PMA_CH0_REG_PLL_READY_OW                 ("DISABLE"                     ),                 
    .PMA_CH0_REG_PLL_READY                    ("TRUE"                        ),                    
    .PMA_CH0_REG_TX_PCLK_SW_OW                ("DISABLE"                     ),                
    .PMA_CH0_REG_TX_PCLK_SW                   ("TRUE"                        ),                   
    .PMA_CH0_REG_EI_PCLK_DELAY_SEL            (0                             ),              
    .PMA_CH0_REG_TX_DRV01_DAC0                (0                             ), 
    .PMA_CH0_REG_TX_DRV01_DAC1                (0                             ), 
    .PMA_CH0_REG_TX_DRV01_DAC2                (0                             ), 
    .PMA_CH0_REG_TX_DRV00_DAC0                (63                            ),                
    .PMA_CH0_REG_TX_DRV00_DAC1                (53                            ),                
    .PMA_CH0_REG_TX_DRV00_DAC2                (48                            ),                
    .PMA_CH0_REG_TX_AMP1                      (16                            ),                      
    .PMA_CH0_REG_TX_AMP2                      (32                            ),                      
    .PMA_CH0_REG_TX_AMP3                      (48                            ),                      
    .PMA_CH0_REG_TX_AMP4                      (56                            ),                      
    .PMA_CH0_REG_TX_MARGIN                    (0                             ),                    
    .PMA_CH0_REG_TX_MARGIN_OW                 ("DISABLE"                     ),                 
    .PMA_CH0_REG_TX_DEEMP                     (0                             ),                     
    .PMA_CH0_REG_TX_DEEMP_OW                  ("DISABLE"                     ),                  
    .PMA_CH0_REG_TX_SWING                     ("FALSE"                       ),                     
    .PMA_CH0_REG_TX_SWING_OW                  ("DISABLE"                     ),                  
    .PMA_CH0_REG_TX_RXDET_THRESHOLD           ("50MV"                        ),           
    .PMA_CH0_REG_TX_BEACON_OSC_CTRL           (4                             ),           
    .PMA_CH0_REG_TX_PREDRV_DAC                (1                             ),                
    .PMA_CH0_REG_TX_PREDRV_CM_CTRL            (1                             ),            
    .PMA_CH0_REG_TX_TX2RX_SLPBACK_EN          ("FALSE"                       ),          
    .PMA_CH0_REG_TX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH0_REG_TX_RXDET_STATUS_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_TX_RXDET_STATUS              ("TRUE"                        ),              
    .PMA_CH0_REG_TX_PRBS_GEN_EN               ("FALSE"                       ),                 
    .PMA_CH0_REG_TX_PRBS_GEN_WIDTH_SEL        ("16BIT"                       ),        
    .PMA_CH0_REG_TX_PRBS_SEL                  ("PRBS7"                       ),                  
    .PMA_CH0_REG_TX_UDP_DATA                  (256773                        ),                  
    .PMA_CH0_REG_TX_FIFO_RST_N                ("FALSE"                       ),                
    .PMA_CH0_REG_TX_FIFO_WP_CTRL              (2                             ),              
    .PMA_CH0_REG_TX_FIFO_EN                   ("FALSE"                       ),                   
    .PMA_CH0_REG_TX_DATA_MUX_SEL              (0                             ),              
    .PMA_CH0_REG_TX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH0_REG_TX_SATA_EN                   ("FALSE"                       ),                   
    .PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON_OW     ("DISABLE"                     ),     
    .PMA_CH0_REG_RATE_CHANGE_TXPCLK_ON        ("ENABLE"                      ),        
    .PMA_CH0_REG_TX_PULLUP_DAC0               (8                             ),               
    .PMA_CH0_REG_TX_PULLUP_DAC1               (8                             ),               
    .PMA_CH0_REG_TX_PULLUP_DAC2               (8                             ),               
    .PMA_CH0_REG_TX_PULLUP_DAC3               (8                             ),               
    .PMA_CH0_REG_TX_OOB_DELAY_SEL             (0                             ),             
    .PMA_CH0_REG_TX_POLARITY                  ("NORMAL"                      ),                  
    .PMA_CH0_REG_TX_SLPBK_AMP                 (1                             ),                 
    .PMA_CH0_REG_TX_LS_MODE_EN                ("FALSE"                       ),                
    .PMA_CH0_REG_TX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_TX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH0_REG_RX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH0_REG_RX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH0_REG_RX_JTAG_OE                   ("DISABLE"                     ),                   
    .PMA_CH0_REG_RX_ACJTAG_VHYSTSE            (0                             ),            
    .PMA_CH0_REG_TX_FBCLK_FAR_EN              ("FALSE"                       ),                
    .PMA_CH0_REG_RX_TERM_MODE_CTRL            (6                             ), 
    .PMA_CH0_REG_PLPBK_TXPCLK_EN              ("TRUE"                        ),              
    .PMA_CH0_REG_TX_609_600                   (0                             ),             
    .PMA_CH0_REG_RX_CDR_617_610               (0                             ),             
    .PMA_CH0_REG_RX_CDR_623_618               (0                             ),             
    .PMA_CH0_REG_RX_631_624                   (0                             ),             
    .PMA_CH0_REG_RX_639_632                   (0                             ),             
    .PMA_CH0_REG_RX_647_640                   (0                             ),             
    .PMA_CH0_REG_RX_655_648                   (0                             ),             
    .PMA_CH0_REG_RX_659_656                   (8                             ),             
    .PMA_CH0_CFG_LANE_POWERUP                 ("ON"                          ),                 
    .PMA_CH0_CFG_PMA_POR_N                    ("TRUE"                        ),                    
    .PMA_CH0_CFG_RX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH0_CFG_RX_PMA_RSTN                  ("TRUE"                        ),                  
    .PMA_CH0_CFG_TX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH0_CFG_TX_PMA_RSTN                  ("TRUE"                        ), 
    .PMA_CH0_CFG_CTLE_ADP_RSTN                ("TRUE"                        ),                 
    .PMA_CH0_REG_RESERVED_48_45               (0                             ),               
    .PMA_CH0_REG_RESERVED_69                  (0                             ),                  
    .PMA_CH0_REG_RESERVED_77_76               (0                             ),               
    .PMA_CH0_REG_RESERVED_171_164             (0                             ),             
    .PMA_CH0_REG_RESERVED_175_172             (0                             ),             
    .PMA_CH0_REG_RESERVED_190                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_233_232             (0                             ),             
    .PMA_CH0_REG_RESERVED_235_234             (0                             ),             
    .PMA_CH0_REG_RESERVED_241_240             (0                             ),             
    .PMA_CH0_REG_RESERVED_285_283             (0                             ),             
    .PMA_CH0_REG_RESERVED_286                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_295                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_298                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_332_325             (0                             ),             
    .PMA_CH0_REG_RESERVED_340_333             (0                             ),             
    .PMA_CH0_REG_RESERVED_348_341             (0                             ),             
    .PMA_CH0_REG_RESERVED_354_349             (0                             ),             
    .PMA_CH0_REG_RESERVED_373                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_376                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_452                 (0                             ),                 
    .PMA_CH0_REG_RESERVED_502_499             (0                             ),             
    .PMA_CH0_REG_RESERVED_506_505             (0                             ),             
    .PMA_CH0_REG_RESERVED_550_549             (0                             ),             
    .PMA_CH0_REG_RESERVED_556_552             (0                             ),             
    .PMA_CH1_REG_RX_PD                        ("ON"                          ),                        
    .PMA_CH1_REG_RX_PD_EN                     ("FALSE"                       ),                     
    .PMA_CH1_REG_RX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH1_REG_RX_CLKPATH_PD_EN             ("FALSE"                       ),             
    .PMA_CH1_REG_RX_DATAPATH_PD               ("ON"                          ),               
    .PMA_CH1_REG_RX_DATAPATH_PD_EN            ("FALSE"                       ),            
    .PMA_CH1_REG_RX_SIGDET_PD                 ("ON"                          ),                 
    .PMA_CH1_REG_RX_SIGDET_PD_EN              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_DCC_RST_N                 ("TRUE"                        ),                 
    .PMA_CH1_REG_RX_DCC_RST_N_EN              ("TRUE"                        ),              
    .PMA_CH1_REG_RX_CDR_RST_N                 ("TRUE"                        ),                 
    .PMA_CH1_REG_RX_CDR_RST_N_EN              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_SIGDET_RST_N              ("TRUE"                        ),              
    .PMA_CH1_REG_RX_SIGDET_RST_N_EN           ("FALSE"                       ),           
    .PMA_CH1_REG_RXPCLK_SLIP                  ("FALSE"                       ),                  
    .PMA_CH1_REG_RXPCLK_SLIP_OW               ("DISABLE"                     ),               
    .PMA_CH1_REG_RX_PCLKSWITCH_RST_N          ("TRUE"                        ),          
    .PMA_CH1_REG_RX_PCLKSWITCH_RST_N_EN       ("FALSE"                       ),       
    .PMA_CH1_REG_RX_PCLKSWITCH                ("FALSE"                       ),                
    .PMA_CH1_REG_RX_PCLKSWITCH_EN             ("FALSE"                       ),               
    .PMA_CH1_REG_RX_HIGHZ                     ("FALSE"                       ), 
    .PMA_CH1_REG_RX_HIGHZ_EN                  ("FALSE"                       ), 
    .PMA_CH1_REG_RX_EQ_C_SET                  (0                             ),                  
    .PMA_CH1_REG_RX_EQ_R_SET                  (1                             ),                    
    .PMA_CH1_REG_RX_BUSWIDTH                  ("16BIT"                       ), 
    .PMA_CH1_REG_RX_BUSWIDTH_EN               ("TRUE"                        ), 
    .PMA_CH1_REG_RX_RATE                      ("DIV4"                        ),                      
    .PMA_CH1_REG_RX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_RX_RES_TRIM                  (51                            ),                  
    .PMA_CH1_REG_RX_RES_TRIM_EN               ("FALSE"                       ),               
    .PMA_CH1_REG_RX_EQ_OFF                    ("FALSE"                       ),                    
    .PMA_CH1_REG_RX_PREAMP_IC                 (1367                          ),                 
    .PMA_CH1_REG_RX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH1_REG_RX_PIBUF_IC                  (2                             ),                  
    .PMA_CH1_REG_RX_DCC_IC_RX                 (3                             ),                 
    .PMA_CH1_REG_RX_DCC_IC_TX                 (3                             ),                 
    .PMA_CH1_REG_RX_ICTRL_TRX                 ("100PCT"                      ),                 
    .PMA_CH1_REG_RX_ICTRL_PREAMP              ("100PCT"                      ),              
    .PMA_CH1_REG_RX_ICTRL_SLICER              ("100PCT"                      ),              
    .PMA_CH1_REG_RX_ICTRL_PIBUF               ("100PCT"                      ),               
    .PMA_CH1_REG_RX_ICTRL_PI                  ("100PCT"                      ),                  
    .PMA_CH1_REG_RX_ICTRL_DCC                 ("100PCT"                      ),                 
    .PMA_CH1_REG_RX_ICTRL_PREDRV              ("100PCT"                      ),                
    .PMA_CH1_REG_TX_RATE                      ("DIV4"                        ),                      
    .PMA_CH1_REG_TX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N         ("TRUE"                        ),         
    .PMA_CH1_REG_RX_TX2RX_PLPBK_RST_N_EN      ("FALSE"                       ),      
    .PMA_CH1_REG_RX_TX2RX_PLPBK_EN            ("FALSE"                       ),            
    .PMA_CH1_REG_TXCLK_SEL                    ("PLL"                         ),                    
    .PMA_CH1_REG_RX_DATA_POLARITY             ("NORMAL"                      ),             
    .PMA_CH1_REG_RX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH1_REG_UDP_CHK_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_PRBS_SEL                     ("PRBS7"                       ),                     
    .PMA_CH1_REG_PRBS_CHK_EN                  ("FALSE"                       ),                     
    .PMA_CH1_REG_PRBS_CHK_WIDTH_SEL           ("16BIT"                       ),            
    .PMA_CH1_REG_BIST_CHK_PAT_SEL             ("PRBS"                        ),             
    .PMA_CH1_REG_LOAD_ERR_CNT                 ("DISABLE"                     ),                 
    .PMA_CH1_REG_CHK_COUNTER_EN               ("FALSE"                       ),               
    .PMA_CH1_REG_CDR_PROP_TURBO_GAIN          (6                             ),          
    .PMA_CH1_REG_CDR_INT_GAIN                 (5                             ),                 
    .PMA_CH1_REG_CDR_INT_TURBO_GAIN           (6                             ),           
    .PMA_CH1_REG_CDR_INT_SAT_MAX              (992                           ),              
    .PMA_CH1_REG_CDR_INT_SAT_MIN              (32                            ),              
    .PMA_CH1_REG_CDR_INT_RST                  ("FALSE"                       ),                  
    .PMA_CH1_REG_CDR_INT_RST_OW               ("DISABLE"                     ),               
    .PMA_CH1_REG_CDR_PROP_RST                 ("FALSE"                       ),                 
    .PMA_CH1_REG_CDR_PROP_RST_OW              ("DISABLE"                     ),              
    .PMA_CH1_REG_CDR_LOCK_RST                 ("FALSE"                       ),                 
    .PMA_CH1_REG_CDR_LOCK_RST_OW              ("DISABLE"                     ),              
    .PMA_CH1_REG_CDR_RX_PI_FORCE_SEL          (0                             ),          
    .PMA_CH1_REG_CDR_RX_PI_FORCE_D            (0                             ),              
    .PMA_CH1_REG_CDR_LOCK_TIMER               ("25_6U"                       ), 
    .PMA_CH1_REG_CDR_TURBO_MODE_TIMER         (1                             ),         
    .PMA_CH1_REG_CDR_LOCK_VAL                 ("FALSE"                       ),                 
    .PMA_CH1_REG_CDR_LOCK_OW                  ("DISABLE"                     ),                  
    .PMA_CH1_REG_CDR_INT_SAT_DET_EN           ("TRUE"                        ),           
    .PMA_CH1_REG_CDR_SAT_DET_STATUS_EN        ("FALSE"                       ),        
    .PMA_CH1_REG_CDR_SAT_DET_STATUS_RESET_EN  ("FALSE"                       ),   
    .PMA_CH1_REG_CDR_PI_CTRL_RST              ("FALSE"                       ),              
    .PMA_CH1_REG_CDR_PI_CTRL_RST_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_CDR_SAT_DET_RST              ("FALSE"                       ),              
    .PMA_CH1_REG_CDR_SAT_DET_RST_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_CDR_SAT_DET_STICKY_RST       ("FALSE"                       ),       
    .PMA_CH1_REG_CDR_SAT_DET_STICKY_RST_OW    ("DISABLE"                     ),    
    .PMA_CH1_REG_CDR_SIGDET_STATUS_DIS        ("FALSE"                       ),        
    .PMA_CH1_REG_CDR_SAT_DET_TIMER            (2                             ),            
    .PMA_CH1_REG_CDR_SAT_DET_STATUS_VAL       ("FALSE"                       ),       
    .PMA_CH1_REG_CDR_SAT_DET_STATUS_OW        ("DISABLE"                     ),        
    .PMA_CH1_REG_CDR_TURBO_MODE_EN            ("TRUE"                        ),            
    .PMA_CH1_REG_CDR_STATUS_RADDR_INIT        (0                             ),        
    .PMA_CH1_REG_CDR_STATUS_FIFO_EN           ("TRUE"                        ),           
    .PMA_CH1_REG_PMA_TEST_SEL                 (0                             ),                 
    .PMA_CH1_REG_OOB_COMWAKE_GAP_MIN          (3                             ),          
    .PMA_CH1_REG_OOB_COMWAKE_GAP_MAX          (11                            ),          
    .PMA_CH1_REG_OOB_COMINIT_GAP_MIN          (15                            ),          
    .PMA_CH1_REG_OOB_COMINIT_GAP_MAX          (35                            ),          
    .PMA_CH1_REG_RX_PIBUF_IC_TX               (1                             ),               
    .PMA_CH1_REG_COMWAKE_STATUS_CLEAR         (0                             ),         
    .PMA_CH1_REG_COMINIT_STATUS_CLEAR         (0                             ),         
    .PMA_CH1_REG_RX_SYNC_RST_N_EN             ("FALSE"                       ),             
    .PMA_CH1_REG_RX_SYNC_RST_N                ("TRUE"                        ),                
    .PMA_CH1_REG_RX_SATA_COMINIT_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_RX_SATA_COMINIT              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_SATA_COMWAKE_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_RX_SATA_COMWAKE              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH1_REG_TX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH1_REG_RX_SLIP_SEL_EN               ("FALSE"                       ),               
    .PMA_CH1_REG_RX_SLIP_SEL                  (0                             ),                  
    .PMA_CH1_REG_RX_SLIP_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_RX_SIGDET_STATUS_SEL         (5                             ),         
    .PMA_CH1_REG_RX_SIGDET_FSM_RST_N          ("TRUE"                        ),          
    .PMA_CH1_REG_RX_SIGDET_STATUS_OW          ("DISABLE"                     ),          
    .PMA_CH1_REG_RX_SIGDET_STATUS             ("FALSE"                       ),             
    .PMA_CH1_REG_RX_SIGDET_GRM                (0                             ),                
    .PMA_CH1_REG_RX_SIGDET_PULSE_EXT          ("DISABLE"                     ),          
    .PMA_CH1_REG_RX_SIGDET_CH2_SEL            (0                             ),            
    .PMA_CH1_REG_RX_SIGDET_CH2_CHK_WINDOW     (3                             ),     
    .PMA_CH1_REG_RX_SIGDET_CHK_WINDOW_EN      ("TRUE"                        ),      
    .PMA_CH1_REG_RX_SIGDET_NOSIG_COUNT_SETTING(4                             ),
    .PMA_CH1_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (0                             ),  
    .PMA_CH1_REG_SLIP_FIFO_INV_EN             ("FALSE"                       ),             
    .PMA_CH1_REG_SLIP_FIFO_INV                ("POS_EDGE"                    ),                
    .PMA_CH1_REG_RX_SIGDET_4OOB_DET_SEL       (7                             ),       
    .PMA_CH1_REG_RX_SIGDET_IC_I               (10                            ),               
    .PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N_OW   ("DISABLE"                     ),   
    .PMA_CH1_REG_RX_OOB_DETECTOR_RESET_N      ("FALSE"                       ),      
    .PMA_CH1_REG_RX_OOB_DETECTOR_PD_OW        ("DISABLE"                     ),        
    .PMA_CH1_REG_RX_OOB_DETECTOR_PD           ("ON"                          ),           
    .PMA_CH1_REG_RX_TERM_CM_CTRL              ("5DIV7"                       ),              
    .PMA_CH1_REG_TX_PD                        ("ON"                          ),                        
    .PMA_CH1_REG_TX_PD_OW                     ("DISABLE"                     ),                     
    .PMA_CH1_REG_TX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH1_REG_TX_CLKPATH_PD_OW             ("DISABLE"                     ),             
    .PMA_CH1_REG_TX_BEACON_TIMER_SEL          (0                             ),          
    .PMA_CH1_REG_TX_RXDET_REQ_OW              ("DISABLE"                     ),              
    .PMA_CH1_REG_TX_RXDET_REQ                 ("FALSE"                       ),                 
    .PMA_CH1_REG_TX_BEACON_EN_OW              ("DISABLE"                     ),              
    .PMA_CH1_REG_TX_BEACON_EN                 ("FALSE"                       ),                 
    .PMA_CH1_REG_TX_EI_EN_OW                  ("DISABLE"                     ),                  
    .PMA_CH1_REG_TX_EI_EN                     ("FALSE"                       ),                     
    .PMA_CH1_REG_TX_RES_CAL_EN                ("FALSE"                       ),                
    .PMA_CH1_REG_TX_RES_CAL                   (51                            ),                   
    .PMA_CH1_REG_TX_BIAS_CAL_EN               ("FALSE"                       ),               
    .PMA_CH1_REG_TX_BIAS_CTRL                 (48                            ),                 
    .PMA_CH1_REG_TX_RXDET_TIMER_SEL           ("12CYCLE"                     ),           
    .PMA_CH1_REG_TX_SYNC_OW                   ("DISABLE"                     ),                   
    .PMA_CH1_REG_TX_SYNC                      ("DISABLE"                     ),                        
    .PMA_CH1_REG_TX_PD_POST                   ("OFF"                         ), 
    .PMA_CH1_REG_TX_PD_POST_OW                ("ENABLE"                      ),               
    .PMA_CH1_REG_TX_RESET_N_OW                ("DISABLE"                     ),                
    .PMA_CH1_REG_TX_RESET_N                   ("TRUE"                        ),                   
    .PMA_CH1_REG_TX_DCC_RESET_N_OW            ("DISABLE"                     ),            
    .PMA_CH1_REG_TX_DCC_RESET_N               ("TRUE"                        ),                 
    .PMA_CH1_REG_TX_BUSWIDTH_OW               ("ENABLE"                      ), 
    .PMA_CH1_REG_TX_BUSWIDTH                  ("16BIT"                       ), 
    .PMA_CH1_REG_PLL_READY_OW                 ("DISABLE"                     ),                 
    .PMA_CH1_REG_PLL_READY                    ("TRUE"                        ),                    
    .PMA_CH1_REG_TX_PCLK_SW_OW                ("DISABLE"                     ),                
    .PMA_CH1_REG_TX_PCLK_SW                   ("TRUE"                        ),                   
    .PMA_CH1_REG_EI_PCLK_DELAY_SEL            (0                             ),              
    .PMA_CH1_REG_TX_DRV01_DAC0                (0                             ), 
    .PMA_CH1_REG_TX_DRV01_DAC1                (0                             ), 
    .PMA_CH1_REG_TX_DRV01_DAC2                (0                             ), 
    .PMA_CH1_REG_TX_DRV00_DAC0                (63                            ),                
    .PMA_CH1_REG_TX_DRV00_DAC1                (53                            ),                
    .PMA_CH1_REG_TX_DRV00_DAC2                (48                            ),                
    .PMA_CH1_REG_TX_AMP1                      (16                            ),                      
    .PMA_CH1_REG_TX_AMP2                      (32                            ),                      
    .PMA_CH1_REG_TX_AMP3                      (48                            ),                      
    .PMA_CH1_REG_TX_AMP4                      (56                            ),                      
    .PMA_CH1_REG_TX_MARGIN                    (0                             ),                    
    .PMA_CH1_REG_TX_MARGIN_OW                 ("DISABLE"                     ),                 
    .PMA_CH1_REG_TX_DEEMP                     (0                             ),                     
    .PMA_CH1_REG_TX_DEEMP_OW                  ("DISABLE"                     ),                  
    .PMA_CH1_REG_TX_SWING                     ("FALSE"                       ),                     
    .PMA_CH1_REG_TX_SWING_OW                  ("DISABLE"                     ),                  
    .PMA_CH1_REG_TX_RXDET_THRESHOLD           ("50MV"                        ),           
    .PMA_CH1_REG_TX_BEACON_OSC_CTRL           (4                             ),           
    .PMA_CH1_REG_TX_PREDRV_DAC                (1                             ),                
    .PMA_CH1_REG_TX_PREDRV_CM_CTRL            (1                             ),            
    .PMA_CH1_REG_TX_TX2RX_SLPBACK_EN          ("FALSE"                       ),          
    .PMA_CH1_REG_TX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH1_REG_TX_RXDET_STATUS_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_TX_RXDET_STATUS              ("TRUE"                        ),              
    .PMA_CH1_REG_TX_PRBS_GEN_EN               ("FALSE"                       ),                 
    .PMA_CH1_REG_TX_PRBS_GEN_WIDTH_SEL        ("16BIT"                       ),          
    .PMA_CH1_REG_TX_PRBS_SEL                  ("PRBS7"                       ),                  
    .PMA_CH1_REG_TX_UDP_DATA                  (256773                        ),                  
    .PMA_CH1_REG_TX_FIFO_RST_N                ("FALSE"                       ),                
    .PMA_CH1_REG_TX_FIFO_WP_CTRL              (2                             ),              
    .PMA_CH1_REG_TX_FIFO_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_TX_DATA_MUX_SEL              (0                             ),              
    .PMA_CH1_REG_TX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH1_REG_TX_SATA_EN                   ("FALSE"                       ),                   
    .PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON_OW     ("DISABLE"                     ),     
    .PMA_CH1_REG_RATE_CHANGE_TXPCLK_ON        ("ENABLE"                      ),        
    .PMA_CH1_REG_TX_PULLUP_DAC0               (8                             ),               
    .PMA_CH1_REG_TX_PULLUP_DAC1               (8                             ),               
    .PMA_CH1_REG_TX_PULLUP_DAC2               (8                             ),               
    .PMA_CH1_REG_TX_PULLUP_DAC3               (8                             ),               
    .PMA_CH1_REG_TX_OOB_DELAY_SEL             (0                             ),             
    .PMA_CH1_REG_TX_POLARITY                  ("NORMAL"                      ),                  
    .PMA_CH1_REG_TX_SLPBK_AMP                 (1                             ),                 
    .PMA_CH1_REG_TX_LS_MODE_EN                ("FALSE"                       ),                
    .PMA_CH1_REG_TX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_TX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH1_REG_RX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH1_REG_RX_JTAG_OE                   ("DISABLE"                     ),                   
    .PMA_CH1_REG_RX_ACJTAG_VHYSTSE            (0                             ),            
    .PMA_CH1_REG_TX_FBCLK_FAR_EN              ("FALSE"                       ),                
    .PMA_CH1_REG_RX_TERM_MODE_CTRL            (6                             ), 
    .PMA_CH1_REG_PLPBK_TXPCLK_EN              ("TRUE"                        ),              
    .PMA_CH1_REG_TX_609_600                   (0                             ),             
    .PMA_CH1_REG_RX_CDR_617_610               (0                             ),             
    .PMA_CH1_REG_RX_CDR_623_618               (0                             ),             
    .PMA_CH1_REG_RX_631_624                   (0                             ),             
    .PMA_CH1_REG_RX_639_632                   (0                             ),             
    .PMA_CH1_REG_RX_647_640                   (0                             ),             
    .PMA_CH1_REG_RX_655_648                   (0                             ),             
    .PMA_CH1_REG_RX_659_656                   (8                             ),             
    .PMA_CH1_CFG_LANE_POWERUP                 ("ON"                          ),                 
    .PMA_CH1_CFG_PMA_POR_N                    ("TRUE"                        ),                    
    .PMA_CH1_CFG_RX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH1_CFG_RX_PMA_RSTN                  ("TRUE"                        ),                  
    .PMA_CH1_CFG_TX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH1_CFG_TX_PMA_RSTN                  ("TRUE"                        ), 
    .PMA_CH1_CFG_CTLE_ADP_RSTN                ("TRUE"                        ),                 
    .PMA_CH1_REG_RESERVED_48_45               (0                             ),               
    .PMA_CH1_REG_RESERVED_69                  (0                             ),                  
    .PMA_CH1_REG_RESERVED_77_76               (0                             ),               
    .PMA_CH1_REG_RESERVED_171_164             (0                             ),             
    .PMA_CH1_REG_RESERVED_175_172             (0                             ),             
    .PMA_CH1_REG_RESERVED_190                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_233_232             (0                             ),             
    .PMA_CH1_REG_RESERVED_235_234             (0                             ),             
    .PMA_CH1_REG_RESERVED_241_240             (0                             ),             
    .PMA_CH1_REG_RESERVED_285_283             (0                             ),             
    .PMA_CH1_REG_RESERVED_286                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_295                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_298                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_332_325             (0                             ),             
    .PMA_CH1_REG_RESERVED_340_333             (0                             ),             
    .PMA_CH1_REG_RESERVED_348_341             (0                             ),             
    .PMA_CH1_REG_RESERVED_354_349             (0                             ),             
    .PMA_CH1_REG_RESERVED_373                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_376                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_452                 (0                             ),                 
    .PMA_CH1_REG_RESERVED_502_499             (0                             ),             
    .PMA_CH1_REG_RESERVED_506_505             (0                             ),             
    .PMA_CH1_REG_RESERVED_550_549             (0                             ),             
    .PMA_CH1_REG_RESERVED_556_552             (0                             ),             
    .PMA_CH2_REG_RX_PD                        ("ON"                          ),                        
    .PMA_CH2_REG_RX_PD_EN                     ("FALSE"                       ),                     
    .PMA_CH2_REG_RX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH2_REG_RX_CLKPATH_PD_EN             ("FALSE"                       ),             
    .PMA_CH2_REG_RX_DATAPATH_PD               ("ON"                          ),               
    .PMA_CH2_REG_RX_DATAPATH_PD_EN            ("FALSE"                       ),            
    .PMA_CH2_REG_RX_SIGDET_PD                 ("ON"                          ),                 
    .PMA_CH2_REG_RX_SIGDET_PD_EN              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_DCC_RST_N                 ("TRUE"                        ),                 
    .PMA_CH2_REG_RX_DCC_RST_N_EN              ("TRUE"                        ),              
    .PMA_CH2_REG_RX_CDR_RST_N                 ("TRUE"                        ),                 
    .PMA_CH2_REG_RX_CDR_RST_N_EN              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_SIGDET_RST_N              ("TRUE"                        ),              
    .PMA_CH2_REG_RX_SIGDET_RST_N_EN           ("FALSE"                       ),           
    .PMA_CH2_REG_RXPCLK_SLIP                  ("FALSE"                       ),                  
    .PMA_CH2_REG_RXPCLK_SLIP_OW               ("DISABLE"                     ),               
    .PMA_CH2_REG_RX_PCLKSWITCH_RST_N          ("TRUE"                        ),          
    .PMA_CH2_REG_RX_PCLKSWITCH_RST_N_EN       ("FALSE"                       ),       
    .PMA_CH2_REG_RX_PCLKSWITCH                ("FALSE"                       ),                
    .PMA_CH2_REG_RX_PCLKSWITCH_EN             ("FALSE"                       ),               
    .PMA_CH2_REG_RX_HIGHZ                     ("FALSE"                       ), 
    .PMA_CH2_REG_RX_HIGHZ_EN                  ("FALSE"                       ), 
    .PMA_CH2_REG_RX_EQ_C_SET                  (0                             ),                  
    .PMA_CH2_REG_RX_EQ_R_SET                  (1                             ),                    
    .PMA_CH2_REG_RX_BUSWIDTH                  ("20BIT"                       ), 
    .PMA_CH2_REG_RX_BUSWIDTH_EN               ("TRUE"                        ), 
    .PMA_CH2_REG_RX_RATE                      ("DIV1"                        ),                      
    .PMA_CH2_REG_RX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH2_REG_RX_RES_TRIM                  (51                            ),                  
    .PMA_CH2_REG_RX_RES_TRIM_EN               ("FALSE"                       ),               
    .PMA_CH2_REG_RX_EQ_OFF                    ("FALSE"                       ),                    
    .PMA_CH2_REG_RX_PREAMP_IC                 (1367                          ),                 
    .PMA_CH2_REG_RX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH2_REG_RX_PIBUF_IC                  (2                             ),                  
    .PMA_CH2_REG_RX_DCC_IC_RX                 (3                             ),                 
    .PMA_CH2_REG_RX_DCC_IC_TX                 (3                             ),                 
    .PMA_CH2_REG_RX_ICTRL_TRX                 ("100PCT"                      ),                 
    .PMA_CH2_REG_RX_ICTRL_PREAMP              ("100PCT"                      ),              
    .PMA_CH2_REG_RX_ICTRL_SLICER              ("100PCT"                      ),              
    .PMA_CH2_REG_RX_ICTRL_PIBUF               ("100PCT"                      ),               
    .PMA_CH2_REG_RX_ICTRL_PI                  ("100PCT"                      ),                  
    .PMA_CH2_REG_RX_ICTRL_DCC                 ("100PCT"                      ),                 
    .PMA_CH2_REG_RX_ICTRL_PREDRV              ("100PCT"                      ),              
    .PMA_CH2_REG_TX_RATE                      ("DIV1"                        ),                      
    .PMA_CH2_REG_TX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N         ("TRUE"                        ),         
    .PMA_CH2_REG_RX_TX2RX_PLPBK_RST_N_EN      ("FALSE"                       ),      
    .PMA_CH2_REG_RX_TX2RX_PLPBK_EN            ("FALSE"                       ),            
    .PMA_CH2_REG_TXCLK_SEL                    ("PLL"                         ),                    
    .PMA_CH2_REG_RX_DATA_POLARITY             ("NORMAL"                      ),             
    .PMA_CH2_REG_RX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH2_REG_UDP_CHK_EN                   ("FALSE"                       ),                   
    .PMA_CH2_REG_PRBS_SEL                     ("PRBS7"                       ),                     
    .PMA_CH2_REG_PRBS_CHK_EN                  ("FALSE"                       ),                   
    .PMA_CH2_REG_PRBS_CHK_WIDTH_SEL           ("20BIT"                       ),          
    .PMA_CH2_REG_BIST_CHK_PAT_SEL             ("PRBS"                        ),             
    .PMA_CH2_REG_LOAD_ERR_CNT                 ("DISABLE"                     ),                 
    .PMA_CH2_REG_CHK_COUNTER_EN               ("FALSE"                       ),               
    .PMA_CH2_REG_CDR_PROP_TURBO_GAIN          (6                             ),          
    .PMA_CH2_REG_CDR_INT_GAIN                 (5                             ),                 
    .PMA_CH2_REG_CDR_INT_TURBO_GAIN           (6                             ),           
    .PMA_CH2_REG_CDR_INT_SAT_MAX              (992                           ),              
    .PMA_CH2_REG_CDR_INT_SAT_MIN              (32                            ),              
    .PMA_CH2_REG_CDR_INT_RST                  ("FALSE"                       ),                  
    .PMA_CH2_REG_CDR_INT_RST_OW               ("DISABLE"                     ),               
    .PMA_CH2_REG_CDR_PROP_RST                 ("FALSE"                       ),                 
    .PMA_CH2_REG_CDR_PROP_RST_OW              ("DISABLE"                     ),              
    .PMA_CH2_REG_CDR_LOCK_RST                 ("FALSE"                       ),                 
    .PMA_CH2_REG_CDR_LOCK_RST_OW              ("DISABLE"                     ),              
    .PMA_CH2_REG_CDR_RX_PI_FORCE_SEL          (0                             ),          
    .PMA_CH2_REG_CDR_RX_PI_FORCE_D            (0                             ),              
    .PMA_CH2_REG_CDR_LOCK_TIMER               ("25_6U"                       ), 
    .PMA_CH2_REG_CDR_TURBO_MODE_TIMER         (1                             ),         
    .PMA_CH2_REG_CDR_LOCK_VAL                 ("FALSE"                       ),                 
    .PMA_CH2_REG_CDR_LOCK_OW                  ("DISABLE"                     ),                  
    .PMA_CH2_REG_CDR_INT_SAT_DET_EN           ("TRUE"                        ),           
    .PMA_CH2_REG_CDR_SAT_DET_STATUS_EN        ("FALSE"                       ),        
    .PMA_CH2_REG_CDR_SAT_DET_STATUS_RESET_EN  ("FALSE"                       ),  
    .PMA_CH2_REG_CDR_PI_CTRL_RST              ("FALSE"                       ),              
    .PMA_CH2_REG_CDR_PI_CTRL_RST_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_CDR_SAT_DET_RST              ("FALSE"                       ),              
    .PMA_CH2_REG_CDR_SAT_DET_RST_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_CDR_SAT_DET_STICKY_RST       ("FALSE"                       ),       
    .PMA_CH2_REG_CDR_SAT_DET_STICKY_RST_OW    ("DISABLE"                     ),    
    .PMA_CH2_REG_CDR_SIGDET_STATUS_DIS        ("FALSE"                       ),        
    .PMA_CH2_REG_CDR_SAT_DET_TIMER            (2                             ),            
    .PMA_CH2_REG_CDR_SAT_DET_STATUS_VAL       ("FALSE"                       ),       
    .PMA_CH2_REG_CDR_SAT_DET_STATUS_OW        ("DISABLE"                     ),        
    .PMA_CH2_REG_CDR_TURBO_MODE_EN            ("TRUE"                        ),            
    .PMA_CH2_REG_CDR_STATUS_RADDR_INIT        (0                             ),        
    .PMA_CH2_REG_CDR_STATUS_FIFO_EN           ("TRUE"                        ),           
    .PMA_CH2_REG_PMA_TEST_SEL                 (0                             ),                 
    .PMA_CH2_REG_OOB_COMWAKE_GAP_MIN          (3                             ),          
    .PMA_CH2_REG_OOB_COMWAKE_GAP_MAX          (11                            ),          
    .PMA_CH2_REG_OOB_COMINIT_GAP_MIN          (15                            ),          
    .PMA_CH2_REG_OOB_COMINIT_GAP_MAX          (35                            ),          
    .PMA_CH2_REG_RX_PIBUF_IC_TX               (1                             ),               
    .PMA_CH2_REG_COMWAKE_STATUS_CLEAR         (0                             ),         
    .PMA_CH2_REG_COMINIT_STATUS_CLEAR         (0                             ),         
    .PMA_CH2_REG_RX_SYNC_RST_N_EN             ("FALSE"                       ),             
    .PMA_CH2_REG_RX_SYNC_RST_N                ("TRUE"                        ),                
    .PMA_CH2_REG_RX_SATA_COMINIT_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_RX_SATA_COMINIT              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_SATA_COMWAKE_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_RX_SATA_COMWAKE              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH2_REG_TX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH2_REG_RX_SLIP_SEL_EN               ("FALSE"                       ),               
    .PMA_CH2_REG_RX_SLIP_SEL                  (0                             ),                  
    .PMA_CH2_REG_RX_SLIP_EN                   ("FALSE"                       ),                   
    .PMA_CH2_REG_RX_SIGDET_STATUS_SEL         (5                             ),         
    .PMA_CH2_REG_RX_SIGDET_FSM_RST_N          ("TRUE"                        ),          
    .PMA_CH2_REG_RX_SIGDET_STATUS_OW          ("DISABLE"                     ),          
    .PMA_CH2_REG_RX_SIGDET_STATUS             ("FALSE"                       ),             
    .PMA_CH2_REG_RX_SIGDET_GRM                (0                             ),                
    .PMA_CH2_REG_RX_SIGDET_PULSE_EXT          ("DISABLE"                     ),          
    .PMA_CH2_REG_RX_SIGDET_CH2_SEL            (0                             ),            
    .PMA_CH2_REG_RX_SIGDET_CH2_CHK_WINDOW     (3                             ),     
    .PMA_CH2_REG_RX_SIGDET_CHK_WINDOW_EN      ("TRUE"                        ),      
    .PMA_CH2_REG_RX_SIGDET_NOSIG_COUNT_SETTING(4                             ),
    .PMA_CH2_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (0                             ),  
    .PMA_CH2_REG_SLIP_FIFO_INV_EN             ("FALSE"                       ),             
    .PMA_CH2_REG_SLIP_FIFO_INV                ("POS_EDGE"                    ),                
    .PMA_CH2_REG_RX_SIGDET_4OOB_DET_SEL       (7                             ),       
    .PMA_CH2_REG_RX_SIGDET_IC_I               (10                            ),               
    .PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N_OW   ("DISABLE"                     ),   
    .PMA_CH2_REG_RX_OOB_DETECTOR_RESET_N      ("FALSE"                       ),      
    .PMA_CH2_REG_RX_OOB_DETECTOR_PD_OW        ("DISABLE"                     ),        
    .PMA_CH2_REG_RX_OOB_DETECTOR_PD           ("ON"                          ),           
    .PMA_CH2_REG_RX_TERM_CM_CTRL              ("5DIV7"                       ),              
    .PMA_CH2_REG_TX_PD                        ("ON"                          ),                        
    .PMA_CH2_REG_TX_PD_OW                     ("DISABLE"                     ),                     
    .PMA_CH2_REG_TX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH2_REG_TX_CLKPATH_PD_OW             ("DISABLE"                     ),             
    .PMA_CH2_REG_TX_BEACON_TIMER_SEL          (0                             ),          
    .PMA_CH2_REG_TX_RXDET_REQ_OW              ("DISABLE"                     ),              
    .PMA_CH2_REG_TX_RXDET_REQ                 ("FALSE"                       ),                 
    .PMA_CH2_REG_TX_BEACON_EN_OW              ("DISABLE"                     ),              
    .PMA_CH2_REG_TX_BEACON_EN                 ("FALSE"                       ),                 
    .PMA_CH2_REG_TX_EI_EN_OW                  ("DISABLE"                     ),                  
    .PMA_CH2_REG_TX_EI_EN                     ("FALSE"                       ),                     
    .PMA_CH2_REG_TX_RES_CAL_EN                ("FALSE"                       ),                
    .PMA_CH2_REG_TX_RES_CAL                   (51                            ),                   
    .PMA_CH2_REG_TX_BIAS_CAL_EN               ("FALSE"                       ),               
    .PMA_CH2_REG_TX_BIAS_CTRL                 (48                            ),                 
    .PMA_CH2_REG_TX_RXDET_TIMER_SEL           ("12CYCLE"                     ),           
    .PMA_CH2_REG_TX_SYNC_OW                   ("DISABLE"                     ),                   
    .PMA_CH2_REG_TX_SYNC                      ("DISABLE"                     ),                        
    .PMA_CH2_REG_TX_PD_POST                   ("OFF"                         ), 
    .PMA_CH2_REG_TX_PD_POST_OW                ("ENABLE"                      ),                
    .PMA_CH2_REG_TX_RESET_N_OW                ("DISABLE"                     ),                
    .PMA_CH2_REG_TX_RESET_N                   ("TRUE"                        ),                   
    .PMA_CH2_REG_TX_DCC_RESET_N_OW            ("DISABLE"                     ),            
    .PMA_CH2_REG_TX_DCC_RESET_N               ("TRUE"                        ),                 
    .PMA_CH2_REG_TX_BUSWIDTH_OW               ("ENABLE"                      ), 
    .PMA_CH2_REG_TX_BUSWIDTH                  ("20BIT"                       ), 
    .PMA_CH2_REG_PLL_READY_OW                 ("DISABLE"                     ),                 
    .PMA_CH2_REG_PLL_READY                    ("TRUE"                        ),                    
    .PMA_CH2_REG_TX_PCLK_SW_OW                ("DISABLE"                     ),                
    .PMA_CH2_REG_TX_PCLK_SW                   ("TRUE"                        ),                   
    .PMA_CH2_REG_EI_PCLK_DELAY_SEL            (0                             ),              
    .PMA_CH2_REG_TX_DRV01_DAC0                (0                             ), 
    .PMA_CH2_REG_TX_DRV01_DAC1                (0                             ), 
    .PMA_CH2_REG_TX_DRV01_DAC2                (0                             ), 
    .PMA_CH2_REG_TX_DRV00_DAC0                (63                            ),                
    .PMA_CH2_REG_TX_DRV00_DAC1                (53                            ),                
    .PMA_CH2_REG_TX_DRV00_DAC2                (48                            ),                
    .PMA_CH2_REG_TX_AMP1                      (16                            ),                      
    .PMA_CH2_REG_TX_AMP2                      (32                            ),                      
    .PMA_CH2_REG_TX_AMP3                      (48                            ),                      
    .PMA_CH2_REG_TX_AMP4                      (56                            ),                      
    .PMA_CH2_REG_TX_MARGIN                    (0                             ),                    
    .PMA_CH2_REG_TX_MARGIN_OW                 ("DISABLE"                     ),                 
    .PMA_CH2_REG_TX_DEEMP                     (0                             ),                     
    .PMA_CH2_REG_TX_DEEMP_OW                  ("DISABLE"                     ),                  
    .PMA_CH2_REG_TX_SWING                     ("FALSE"                       ),                     
    .PMA_CH2_REG_TX_SWING_OW                  ("DISABLE"                     ),                  
    .PMA_CH2_REG_TX_RXDET_THRESHOLD           ("50MV"                        ),           
    .PMA_CH2_REG_TX_BEACON_OSC_CTRL           (4                             ),           
    .PMA_CH2_REG_TX_PREDRV_DAC                (1                             ),                
    .PMA_CH2_REG_TX_PREDRV_CM_CTRL            (1                             ),            
    .PMA_CH2_REG_TX_TX2RX_SLPBACK_EN          ("FALSE"                       ),          
    .PMA_CH2_REG_TX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH2_REG_TX_RXDET_STATUS_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_TX_RXDET_STATUS              ("TRUE"                        ),              
    .PMA_CH2_REG_TX_PRBS_GEN_EN               ("FALSE"                       ),               
    .PMA_CH2_REG_TX_PRBS_GEN_WIDTH_SEL        ("20BIT"                       ),         
    .PMA_CH2_REG_TX_PRBS_SEL                  ("PRBS7"                       ),                  
    .PMA_CH2_REG_TX_UDP_DATA                  (256773                        ),                  
    .PMA_CH2_REG_TX_FIFO_RST_N                ("FALSE"                       ),                
    .PMA_CH2_REG_TX_FIFO_WP_CTRL              (2                             ),              
    .PMA_CH2_REG_TX_FIFO_EN                   ("FALSE"                       ),                   
    .PMA_CH2_REG_TX_DATA_MUX_SEL              (0                             ),              
    .PMA_CH2_REG_TX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH2_REG_TX_SATA_EN                   ("FALSE"                       ),                             
    .PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON_OW     ("DISABLE"                     ),     
    .PMA_CH2_REG_RATE_CHANGE_TXPCLK_ON        ("ENABLE"                      ),        
    .PMA_CH2_REG_TX_PULLUP_DAC0               (8                             ),               
    .PMA_CH2_REG_TX_PULLUP_DAC1               (8                             ),               
    .PMA_CH2_REG_TX_PULLUP_DAC2               (8                             ),               
    .PMA_CH2_REG_TX_PULLUP_DAC3               (8                             ),               
    .PMA_CH2_REG_TX_OOB_DELAY_SEL             (0                             ),             
    .PMA_CH2_REG_TX_POLARITY                  ("NORMAL"                      ),                  
    .PMA_CH2_REG_TX_SLPBK_AMP                 (1                             ),                 
    .PMA_CH2_REG_TX_LS_MODE_EN                ("FALSE"                       ),                
    .PMA_CH2_REG_TX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_TX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_JTAG_MODE_EN_OW           ("DISABLE"                     ),           
    .PMA_CH2_REG_RX_JTAG_MODE_EN              ("FALSE"                       ),              
    .PMA_CH2_REG_RX_JTAG_OE                   ("DISABLE"                     ),                   
    .PMA_CH2_REG_RX_ACJTAG_VHYSTSE            (0                             ),            
    .PMA_CH2_REG_TX_FBCLK_FAR_EN              ("FALSE"                       ),                
    .PMA_CH2_REG_RX_TERM_MODE_CTRL            (6                             ), 
    .PMA_CH2_REG_PLPBK_TXPCLK_EN              ("TRUE"                        ),              
    .PMA_CH2_REG_TX_609_600                   (0                             ),             
    .PMA_CH2_REG_RX_CDR_617_610               (0                             ),             
    .PMA_CH2_REG_RX_CDR_623_618               (0                             ),             
    .PMA_CH2_REG_RX_631_624                   (0                             ),             
    .PMA_CH2_REG_RX_639_632                   (0                             ),             
    .PMA_CH2_REG_RX_647_640                   (0                             ),             
    .PMA_CH2_REG_RX_655_648                   (0                             ),             
    .PMA_CH2_REG_RX_659_656                   (8                             ),             
    .PMA_CH2_CFG_LANE_POWERUP                 ("ON"                          ),                 
    .PMA_CH2_CFG_PMA_POR_N                    ("TRUE"                        ),                    
    .PMA_CH2_CFG_RX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH2_CFG_RX_PMA_RSTN                  ("TRUE"                        ),                  
    .PMA_CH2_CFG_TX_LANE_POWERUP              ("ON"                          ),              
    .PMA_CH2_CFG_TX_PMA_RSTN                  ("TRUE"                        ),                  
    .PMA_CH2_CFG_CTLE_ADP_RSTN                ("TRUE"                        ),
    .PMA_CH2_REG_RESERVED_48_45               (0                             ),               
    .PMA_CH2_REG_RESERVED_69                  (0                             ),                  
    .PMA_CH2_REG_RESERVED_77_76               (0                             ),               
    .PMA_CH2_REG_RESERVED_171_164             (0                             ),             
    .PMA_CH2_REG_RESERVED_175_172             (0                             ),             
    .PMA_CH2_REG_RESERVED_190                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_233_232             (0                             ),             
    .PMA_CH2_REG_RESERVED_235_234             (0                             ),             
    .PMA_CH2_REG_RESERVED_241_240             (0                             ),             
    .PMA_CH2_REG_RESERVED_285_283             (0                             ),             
    .PMA_CH2_REG_RESERVED_286                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_295                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_298                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_332_325             (0                             ),             
    .PMA_CH2_REG_RESERVED_340_333             (0                             ),             
    .PMA_CH2_REG_RESERVED_348_341             (0                             ),             
    .PMA_CH2_REG_RESERVED_354_349             (0                             ),             
    .PMA_CH2_REG_RESERVED_373                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_376                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_452                 (0                             ),                 
    .PMA_CH2_REG_RESERVED_502_499             (0                             ),             
    .PMA_CH2_REG_RESERVED_506_505             (0                             ),             
    .PMA_CH2_REG_RESERVED_550_549             (0                             ),             
    .PMA_CH2_REG_RESERVED_556_552             (0                             ),             
    .PMA_CH3_REG_RX_PD                        ("ON"                          ),                        
    .PMA_CH3_REG_RX_PD_EN                     ("FALSE"                       ),                     
    .PMA_CH3_REG_RX_CLKPATH_PD                ("ON"                          ),                
    .PMA_CH3_REG_RX_CLKPATH_PD_EN             ("FALSE"                       ),             
    .PMA_CH3_REG_RX_DATAPATH_PD               ("ON"                          ),               
    .PMA_CH3_REG_RX_DATAPATH_PD_EN            ("FALSE"                       ),            
    .PMA_CH3_REG_RX_SIGDET_PD                 ("ON"                          ),                 
    .PMA_CH3_REG_RX_SIGDET_PD_EN              ("FALSE"                       ),              
    .PMA_CH3_REG_RX_DCC_RST_N                 ("TRUE"                        ),                 
    .PMA_CH3_REG_RX_DCC_RST_N_EN              ("TRUE"                        ),              
    .PMA_CH3_REG_RX_CDR_RST_N                 ("TRUE"                        ),                 
    .PMA_CH3_REG_RX_CDR_RST_N_EN              ("FALSE"                       ),              
    .PMA_CH3_REG_RX_SIGDET_RST_N              ("TRUE"                        ),              
    .PMA_CH3_REG_RX_SIGDET_RST_N_EN           ("FALSE"                       ),           
    .PMA_CH3_REG_RXPCLK_SLIP                  ("FALSE"                       ),                  
    .PMA_CH3_REG_RXPCLK_SLIP_OW               ("DISABLE"                     ),               
    .PMA_CH3_REG_RX_PCLKSWITCH_RST_N          ("TRUE"                        ),          
    .PMA_CH3_REG_RX_PCLKSWITCH_RST_N_EN       ("FALSE"                       ),       
    .PMA_CH3_REG_RX_PCLKSWITCH                ("FALSE"                       ),                
    .PMA_CH3_REG_RX_PCLKSWITCH_EN             ("FALSE"                       ),               
    .PMA_CH3_REG_RX_HIGHZ                     ("FALSE"                       ), 
    .PMA_CH3_REG_RX_HIGHZ_EN                  ("FALSE"                       ), 
    .PMA_CH3_REG_RX_EQ_C_SET                  (0                             ),                  
    .PMA_CH3_REG_RX_EQ_R_SET                  (1                             ),                    
    .PMA_CH3_REG_RX_BUSWIDTH                  ("20BIT"                       ), 
    .PMA_CH3_REG_RX_BUSWIDTH_EN               ("TRUE"                        ), 
    .PMA_CH3_REG_RX_RATE                      ("DIV1"                        ),                      
    .PMA_CH3_REG_RX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH3_REG_RX_RES_TRIM                  (51                            ),                  
    .PMA_CH3_REG_RX_RES_TRIM_EN               ("FALSE"                       ),               
    .PMA_CH3_REG_RX_EQ_OFF                    ("FALSE"                       ),                    
    .PMA_CH3_REG_RX_PREAMP_IC                 (1367                          ),                 
    .PMA_CH3_REG_RX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),             
    .PMA_CH3_REG_RX_PIBUF_IC                  (2                             ),                  
    .PMA_CH3_REG_RX_DCC_IC_RX                 (3                             ),                 
    .PMA_CH3_REG_RX_DCC_IC_TX                 (3                             ),                 
    .PMA_CH3_REG_RX_ICTRL_TRX                 ("100PCT"                      ),                 
    .PMA_CH3_REG_RX_ICTRL_PREAMP              ("100PCT"                      ),              
    .PMA_CH3_REG_RX_ICTRL_SLICER              ("100PCT"                      ),              
    .PMA_CH3_REG_RX_ICTRL_PIBUF               ("100PCT"                      ),               
    .PMA_CH3_REG_RX_ICTRL_PI                  ("100PCT"                      ),                  
    .PMA_CH3_REG_RX_ICTRL_DCC                 ("100PCT"                      ),                 
    .PMA_CH3_REG_RX_ICTRL_PREDRV              ("100PCT"                      ),              
    .PMA_CH3_REG_TX_RATE                      ("DIV1"                        ),                      
    .PMA_CH3_REG_TX_RATE_EN                   ("FALSE"                       ),                   
    .PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N         ("TRUE"                        ),         
    .PMA_CH3_REG_RX_TX2RX_PLPBK_RST_N_EN      ("FALSE"                       ),      
    .PMA_CH3_REG_RX_TX2RX_PLPBK_EN            ("FALSE"                       ),            
    .PMA_CH3_REG_TXCLK_SEL                    ("PLL"                         ),                    
    .PMA_CH3_REG_RX_DATA_POLARITY             ("NORMAL"                      ),             
    .PMA_CH3_REG_RX_ERR_INSERT                ("FALSE"                       ),                
    .PMA_CH3_REG_UDP_CHK_EN                   ("FALSE"                       ),                   
    .PMA_CH3_REG_PRBS_SEL                     ("PRBS7"                       ),                     
    .PMA_CH3_REG_PRBS_CHK_EN                  ("FALSE"                       ),                 
    .PMA_CH3_REG_PRBS_CHK_WIDTH_SEL           ("20BIT"                       ),           
    .PMA_CH3_REG_BIST_CHK_PAT_SEL             ("PRBS"                        ),             
    .PMA_CH3_REG_LOAD_ERR_CNT                 ("DISABLE"                     ),                 
    .PMA_CH3_REG_CHK_COUNTER_EN               ("FALSE"                       ),               
    .PMA_CH3_REG_CDR_PROP_TURBO_GAIN          (6                             ),          
    .PMA_CH3_REG_CDR_INT_GAIN                 (5                             ),                 
    .PMA_CH3_REG_CDR_INT_TURBO_GAIN           (6                             ),           
    .PMA_CH3_REG_CDR_INT_SAT_MAX              (992                           ),              
    .PMA_CH3_REG_CDR_INT_SAT_MIN              (32                            ),              
    .PMA_CH3_REG_CDR_INT_RST                  ("FALSE"                       ),                  
    .PMA_CH3_REG_CDR_INT_RST_OW               ("DISABLE"                     ),               
    .PMA_CH3_REG_CDR_PROP_RST                 ("FALSE"                       ),                 
    .PMA_CH3_REG_CDR_PROP_RST_OW              ("DISABLE"                     ),              
    .PMA_CH3_REG_CDR_LOCK_RST                 ("FALSE"                       ),                 
    .PMA_CH3_REG_CDR_LOCK_RST_OW              ("DISABLE"                     ),              
    .PMA_CH3_REG_CDR_RX_PI_FORCE_SEL          (0                             ),          
    .PMA_CH3_REG_CDR_RX_PI_FORCE_D            (0                             ),              
    .PMA_CH3_REG_CDR_LOCK_TIMER               ("25_6U"                       ), 
    .PMA_CH3_REG_CDR_TURBO_MODE_TIMER         (1                             ),         
    .PMA_CH3_REG_CDR_LOCK_VAL                 ("FALSE"                       ),                 
    .PMA_CH3_REG_CDR_LOCK_OW                  ("DISABLE"                     ),                  
    .PMA_CH3_REG_CDR_INT_SAT_DET_EN           ("TRUE"                        ),           
    .PMA_CH3_REG_CDR_SAT_DET_STATUS_EN        ("FALSE"                       ),        
    .PMA_CH3_REG_CDR_SAT_DET_STATUS_RESET_EN  ("FALSE"                       ),  
    .PMA_CH3_REG_CDR_PI_CTRL_RST              ("FALSE"                       ),              
    .PMA_CH3_REG_CDR_PI_CTRL_RST_OW           ("DISABLE"                     ),           
    .PMA_CH3_REG_CDR_SAT_DET_RST              ("FALSE"                       ),              
    .PMA_CH3_REG_CDR_SAT_DET_RST_OW           ("DISABLE"                     ),           
    .PMA_CH3_REG_CDR_SAT_DET_STICKY_RST       ("FALSE"                       ),       
    .PMA_CH3_REG_CDR_SAT_DET_STICKY_RST_OW    ("DISABLE"                     ),    
    .PMA_CH3_REG_CDR_SIGDET_STATUS_DIS        ("FALSE"                       ),        
    .PMA_CH3_REG_CDR_SAT_DET_TIMER            (2                             ),            
    .PMA_CH3_REG_CDR_SAT_DET_STATUS_VAL       ("FALSE"                       ),       
    .PMA_CH3_REG_CDR_SAT_DET_STATUS_OW        ("DISABLE"                     ),       
    .PMA_CH3_REG_CDR_TURBO_MODE_EN            ("TRUE"                        ),            
    .PMA_CH3_REG_CDR_STATUS_RADDR_INIT        (0                             ),        
    .PMA_CH3_REG_CDR_STATUS_FIFO_EN           ("TRUE"                        ),           
    .PMA_CH3_REG_PMA_TEST_SEL                 (0                             ),                 
    .PMA_CH3_REG_OOB_COMWAKE_GAP_MIN          (3                             ),          
    .PMA_CH3_REG_OOB_COMWAKE_GAP_MAX          (11                            ),          
    .PMA_CH3_REG_OOB_COMINIT_GAP_MIN          (15                            ),          
    .PMA_CH3_REG_OOB_COMINIT_GAP_MAX          (35                            ),          
    .PMA_CH3_REG_RX_PIBUF_IC_TX               (1                             ),               
    .PMA_CH3_REG_COMWAKE_STATUS_CLEAR         (0                             ),         
    .PMA_CH3_REG_COMINIT_STATUS_CLEAR         (0                             ),         
    .PMA_CH3_REG_RX_SYNC_RST_N_EN             ("FALSE"                       ),             
    .PMA_CH3_REG_RX_SYNC_RST_N                ("TRUE"                        ),                
    .PMA_CH3_REG_RX_SATA_COMINIT_OW           ("DISABLE"                     ),           
    .PMA_CH3_REG_RX_SATA_COMINIT              ("FALSE"                       ),              
    .PMA_CH3_REG_RX_SATA_COMWAKE_OW           ("DISABLE"                     ),           
    .PMA_CH3_REG_RX_SATA_COMWAKE              ("FALSE"                       ),              
    .PMA_CH3_REG_RX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH3_REG_TX_DCC_DISABLE               ("ENABLE"                      ),               
    .PMA_CH3_REG_RX_SLIP_SEL_EN               ("FALSE"                       ),               
    .PMA_CH3_REG_RX_SLIP_SEL                  (0                             ),                  
    .PMA_CH3_REG_RX_SLIP_EN                   ("FALSE"                       ),                   
    .PMA_CH3_REG_RX_SIGDET_STATUS_SEL         (5                             ),         
    .PMA_CH3_REG_RX_SIGDET_FSM_RST_N          ("TRUE"                        ),          
    .PMA_CH3_REG_RX_SIGDET_STATUS_OW          ("DISABLE"                     ),          
    .PMA_CH3_REG_RX_SIGDET_STATUS             ("FALSE"                       ),             
    .PMA_CH3_REG_RX_SIGDET_GRM                (0                             ),                
    .PMA_CH3_REG_RX_SIGDET_PULSE_EXT          ("DISABLE"                     ),          
    .PMA_CH3_REG_RX_SIGDET_CH2_SEL            (0                             ),            
    .PMA_CH3_REG_RX_SIGDET_CH2_CHK_WINDOW     (3                             ),     
    .PMA_CH3_REG_RX_SIGDET_CHK_WINDOW_EN      ("TRUE"                        ),      
    .PMA_CH3_REG_RX_SIGDET_NOSIG_COUNT_SETTING(4                             ),
    .PMA_CH3_REG_RX_SIGDET_OOB_DET_COUNT_VAL  (0                             ),
    .PMA_CH3_REG_SLIP_FIFO_INV_EN             ("FALSE"                       ),          
    .PMA_CH3_REG_SLIP_FIFO_INV                ("POS_EDGE"                    ),             
    .PMA_CH3_REG_RX_SIGDET_4OOB_DET_SEL       (7                             ),    
    .PMA_CH3_REG_RX_SIGDET_IC_I               (10                            ),            
    .PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N_OW   ("DISABLE"                     ),
    .PMA_CH3_REG_RX_OOB_DETECTOR_RESET_N      ("FALSE"                       ),   
    .PMA_CH3_REG_RX_OOB_DETECTOR_PD_OW        ("DISABLE"                     ),     
    .PMA_CH3_REG_RX_OOB_DETECTOR_PD           ("ON"                          ),        
    .PMA_CH3_REG_RX_TERM_CM_CTRL              ("5DIV7"                       ),           
    .PMA_CH3_REG_TX_PD                        ("ON"                          ),                     
    .PMA_CH3_REG_TX_PD_OW                     ("DISABLE"                     ),                  
    .PMA_CH3_REG_TX_CLKPATH_PD                ("ON"                          ),             
    .PMA_CH3_REG_TX_CLKPATH_PD_OW             ("DISABLE"                     ),          
    .PMA_CH3_REG_TX_BEACON_TIMER_SEL          (0                             ),       
    .PMA_CH3_REG_TX_RXDET_REQ_OW              ("DISABLE"                     ),           
    .PMA_CH3_REG_TX_RXDET_REQ                 ("FALSE"                       ),              
    .PMA_CH3_REG_TX_BEACON_EN_OW              ("DISABLE"                     ),           
    .PMA_CH3_REG_TX_BEACON_EN                 ("FALSE"                       ),              
    .PMA_CH3_REG_TX_EI_EN_OW                  ("DISABLE"                     ),               
    .PMA_CH3_REG_TX_EI_EN                     ("FALSE"                       ),                  
    .PMA_CH3_REG_TX_RES_CAL_EN                ("FALSE"                       ),             
    .PMA_CH3_REG_TX_RES_CAL                   (51                            ),                
    .PMA_CH3_REG_TX_BIAS_CAL_EN               ("FALSE"                       ),            
    .PMA_CH3_REG_TX_BIAS_CTRL                 (48                            ),              
    .PMA_CH3_REG_TX_RXDET_TIMER_SEL           ("12CYCLE"                     ),        
    .PMA_CH3_REG_TX_SYNC_OW                   ("DISABLE"                     ),                
    .PMA_CH3_REG_TX_SYNC                      ("DISABLE"                     ),                     
    .PMA_CH3_REG_TX_PD_POST                   ("OFF"                         ), 
    .PMA_CH3_REG_TX_PD_POST_OW                ("ENABLE"                      ),             
    .PMA_CH3_REG_TX_RESET_N_OW                ("DISABLE"                     ),             
    .PMA_CH3_REG_TX_RESET_N                   ("TRUE"                        ),                
    .PMA_CH3_REG_TX_DCC_RESET_N_OW            ("DISABLE"                     ),         
    .PMA_CH3_REG_TX_DCC_RESET_N               ("TRUE"                        ),              
    .PMA_CH3_REG_TX_BUSWIDTH_OW               ("ENABLE"                      ), 
    .PMA_CH3_REG_TX_BUSWIDTH                  ("20BIT"                       ), 
    .PMA_CH3_REG_PLL_READY_OW                 ("DISABLE"                     ),              
    .PMA_CH3_REG_PLL_READY                    ("TRUE"                        ),                 
    .PMA_CH3_REG_TX_PCLK_SW_OW                ("DISABLE"                     ),             
    .PMA_CH3_REG_TX_PCLK_SW                   ("TRUE"                        ),                
    .PMA_CH3_REG_EI_PCLK_DELAY_SEL            (0                             ),           
    .PMA_CH3_REG_TX_DRV01_DAC0                (0                             ), 
    .PMA_CH3_REG_TX_DRV01_DAC1                (0                             ), 
    .PMA_CH3_REG_TX_DRV01_DAC2                (0                             ), 
    .PMA_CH3_REG_TX_DRV00_DAC0                (63                            ),             
    .PMA_CH3_REG_TX_DRV00_DAC1                (53                            ),             
    .PMA_CH3_REG_TX_DRV00_DAC2                (48                            ),             
    .PMA_CH3_REG_TX_AMP1                      (16                            ),                   
    .PMA_CH3_REG_TX_AMP2                      (32                            ),                   
    .PMA_CH3_REG_TX_AMP3                      (48                            ),                   
    .PMA_CH3_REG_TX_AMP4                      (56                            ),                   
    .PMA_CH3_REG_TX_MARGIN                    (0                             ),                 
    .PMA_CH3_REG_TX_MARGIN_OW                 ("DISABLE"                     ),              
    .PMA_CH3_REG_TX_DEEMP                     (0                             ),                  
    .PMA_CH3_REG_TX_DEEMP_OW                  ("DISABLE"                     ),               
    .PMA_CH3_REG_TX_SWING                     ("FALSE"                       ),                  
    .PMA_CH3_REG_TX_SWING_OW                  ("DISABLE"                     ),               
    .PMA_CH3_REG_TX_RXDET_THRESHOLD           ("50MV"                        ),        
    .PMA_CH3_REG_TX_BEACON_OSC_CTRL           (4                             ),        
    .PMA_CH3_REG_TX_PREDRV_DAC                (1                             ),             
    .PMA_CH3_REG_TX_PREDRV_CM_CTRL            (1                             ),         
    .PMA_CH3_REG_TX_TX2RX_SLPBACK_EN          ("FALSE"                       ),       
    .PMA_CH3_REG_TX_PCLK_EDGE_SEL             ("POS_EDGE"                    ),          
    .PMA_CH3_REG_TX_RXDET_STATUS_OW           ("DISABLE"                     ),        
    .PMA_CH3_REG_TX_RXDET_STATUS              ("TRUE"                        ),           
    .PMA_CH3_REG_TX_PRBS_GEN_EN               ("FALSE"                       ),              
    .PMA_CH3_REG_TX_PRBS_GEN_WIDTH_SEL        ("20BIT"                       ),     
    .PMA_CH3_REG_TX_PRBS_SEL                  ("PRBS7"                       ),               
    .PMA_CH3_REG_TX_UDP_DATA                  (256773                        ),               
    .PMA_CH3_REG_TX_FIFO_RST_N                ("FALSE"                       ),             
    .PMA_CH3_REG_TX_FIFO_WP_CTRL              (2                             ),           
    .PMA_CH3_REG_TX_FIFO_EN                   ("FALSE"                       ),                
    .PMA_CH3_REG_TX_DATA_MUX_SEL              (0                             ),           
    .PMA_CH3_REG_TX_ERR_INSERT                ("FALSE"                       ),             
    .PMA_CH3_REG_TX_SATA_EN                   ("FALSE"                       ),                
    .PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON_OW     ("DISABLE"                     ),  
    .PMA_CH3_REG_RATE_CHANGE_TXPCLK_ON        ("ENABLE"                      ),     
    .PMA_CH3_REG_TX_PULLUP_DAC0               (8                             ),            
    .PMA_CH3_REG_TX_PULLUP_DAC1               (8                             ),            
    .PMA_CH3_REG_TX_PULLUP_DAC2               (8                             ),            
    .PMA_CH3_REG_TX_PULLUP_DAC3               (8                             ),            
    .PMA_CH3_REG_TX_OOB_DELAY_SEL             (0                             ),          
    .PMA_CH3_REG_TX_POLARITY                  ("NORMAL"                      ),               
    .PMA_CH3_REG_TX_SLPBK_AMP                 (1                             ),              
    .PMA_CH3_REG_TX_LS_MODE_EN                ("FALSE"                       ),             
    .PMA_CH3_REG_TX_JTAG_MODE_EN_OW           ("DISABLE"                     ),        
    .PMA_CH3_REG_TX_JTAG_MODE_EN              ("FALSE"                       ),           
    .PMA_CH3_REG_RX_JTAG_MODE_EN_OW           ("DISABLE"                     ),        
    .PMA_CH3_REG_RX_JTAG_MODE_EN              ("FALSE"                       ),           
    .PMA_CH3_REG_RX_JTAG_OE                   ("DISABLE"                     ),                
    .PMA_CH3_REG_RX_ACJTAG_VHYSTSE            (0                             ),         
    .PMA_CH3_REG_TX_FBCLK_FAR_EN              ("FALSE"                       ),             
    .PMA_CH3_REG_RX_TERM_MODE_CTRL            (6                             ), 
    .PMA_CH3_REG_PLPBK_TXPCLK_EN              ("TRUE"                        ),           
    .PMA_CH3_REG_TX_609_600                   (0                             ),             
    .PMA_CH3_REG_RX_CDR_617_610               (0                             ),             
    .PMA_CH3_REG_RX_CDR_623_618               (0                             ),             
    .PMA_CH3_REG_RX_631_624                   (0                             ),             
    .PMA_CH3_REG_RX_639_632                   (0                             ),             
    .PMA_CH3_REG_RX_647_640                   (0                             ),             
    .PMA_CH3_REG_RX_655_648                   (0                             ),             
    .PMA_CH3_REG_RX_659_656                   (8                             ),             
    .PMA_CH3_CFG_LANE_POWERUP                 ("ON"                          ),              
    .PMA_CH3_CFG_PMA_POR_N                    ("TRUE"                        ),                 
    .PMA_CH3_CFG_RX_LANE_POWERUP              ("ON"                          ),           
    .PMA_CH3_CFG_RX_PMA_RSTN                  ("TRUE"                        ),               
    .PMA_CH3_CFG_TX_LANE_POWERUP              ("ON"                          ),           
    .PMA_CH3_CFG_CTLE_ADP_RSTN                ("TRUE"                        ),
    .PMA_CH3_CFG_TX_PMA_RSTN                  ("TRUE"                        ),               
    .PMA_CH3_REG_RESERVED_48_45               (0                             ),            
    .PMA_CH3_REG_RESERVED_69                  (0                             ),               
    .PMA_CH3_REG_RESERVED_77_76               (0                             ),            
    .PMA_CH3_REG_RESERVED_171_164             (0                             ),          
    .PMA_CH3_REG_RESERVED_175_172             (0                             ),          
    .PMA_CH3_REG_RESERVED_190                 (0                             ),              
    .PMA_CH3_REG_RESERVED_233_232             (0                             ),          
    .PMA_CH3_REG_RESERVED_235_234             (0                             ),          
    .PMA_CH3_REG_RESERVED_241_240             (0                             ),          
    .PMA_CH3_REG_RESERVED_285_283             (0                             ),          
    .PMA_CH3_REG_RESERVED_286                 (0                             ),              
    .PMA_CH3_REG_RESERVED_295                 (0                             ),              
    .PMA_CH3_REG_RESERVED_298                 (0                             ),              
    .PMA_CH3_REG_RESERVED_332_325             (0                             ),          
    .PMA_CH3_REG_RESERVED_340_333             (0                             ),          
    .PMA_CH3_REG_RESERVED_348_341             (0                             ),          
    .PMA_CH3_REG_RESERVED_354_349             (0                             ),          
    .PMA_CH3_REG_RESERVED_373                 (0                             ),              
    .PMA_CH3_REG_RESERVED_376                 (0                             ),              
    .PMA_CH3_REG_RESERVED_452                 (0                             ),              
    .PMA_CH3_REG_RESERVED_502_499             (0                             ),          
    .PMA_CH3_REG_RESERVED_506_505             (0                             ),          
    .PMA_CH3_REG_RESERVED_550_549             (0                             ),          
    .PMA_CH3_REG_RESERVED_556_552             (0                             ),          
    .PMA_PLL0_REG_PLL_POWERDOWN_OW            ("DISABLE"                     ),         
    .PMA_PLL0_REG_PLL_POWERDOWN               ("ON"                          ),            
    .PMA_PLL0_REG_PLL_RESET_N_OW              ("DISABLE"                     ),           
    .PMA_PLL0_REG_PLL_RESET_N                 ("TRUE"                        ),              
    .PMA_PLL0_REG_PLL_READY_OW                ("DISABLE"                     ),             
    .PMA_PLL0_REG_PLL_READY                   ("FALSE"                       ),                
    .PMA_PLL0_REG_LANE_SYNC_OW                ("DISABLE"                     ),             
    .PMA_PLL0_REG_LANE_SYNC                   ("FALSE"                       ),                
    .PMA_PLL0_REG_LOCKDET_REPEAT              ("DISABLE"                     ),           
    .PMA_PLL0_REG_RESCAL_I_CODE_PMA           ("DISABLE"                     ),        
    .PMA_PLL0_REG_RESCAL_RESET_N_OW           ("DISABLE"                     ),        
    .PMA_PLL0_REG_RESCAL_RESET_N              ("FALSE"                       ),           
    .PMA_PLL0_REG_RESCAL_DONE_OW              ("DISABLE"                     ),           
    .PMA_PLL0_REG_RESCAL_DONE                 ("FALSE"                       ),              
    .PMA_PLL0_REG_RESCAL_CODE_OW              ("DISABLE"                     ),           
    .PMA_PLL0_REG_LDO_VREF_SEL                (2                             ),             
    .PMA_PLL0_REG_BIAS_VCOREP_C               (1                             ),            
    .PMA_PLL0_REG_RESCAL_I_CODE               (32                            ),            
    .PMA_PLL0_REG_RESCAL_ONCHIP_SMALL_OW      ("DISABLE"                     ),   
    .PMA_PLL0_REG_RESCAL_ONCHIP_SMALL         (0                             ),      
    .PMA_PLL0_REG_JTAG_OE                     ("DISABLE"                     ),                  
    .PMA_PLL0_REG_JTAG_AC_MODE                ("DISABLE"                     ),             
    .PMA_PLL0_REG_JTAG_VHYSTSEL               (0                             ),            
    .PMA_PLL0_REG_PLL_LOCKDET_EN_OW           ("DISABLE"                     ),        
    .PMA_PLL0_REG_PLL_LOCKDET_EN              ("FALSE"                       ),           
    .PMA_PLL0_REG_PLL_LOCKDET_RESET_N_OW      ("DISABLE"                     ),   
    .PMA_PLL0_REG_PLL_LOCKDET_RESET_N         ("FALSE"                       ),      
    .PMA_PLL0_REG_PLL_LOCKED_OW               ("DISABLE"                     ),            
    .PMA_PLL0_REG_PLL_LOCKED                  ("FALSE"                       ),               
    .PMA_PLL0_REG_PLL_LOCKED_STICKY_CLEAR     ("FALSE"                       ),  
    .PMA_PLL0_REG_PLL_UNLOCKED_STICKY_CLEAR   ("FALSE"                       ),
    .PMA_PLL0_REG_NOFBCLK_STICKY_CLEAR        ("FALSE"                       ), 
    `ifdef IPML_HSST_SPEEDUP_SIM
    .PMA_PLL0_REG_PLL_LOCKDET_REFCT           (4                             ), 
    .PMA_PLL0_REG_PLL_LOCKDET_FBCT            (4                             ), 
    .PMA_PLL0_REG_PLL_LOCKDET_ITER            (0                             ),
    `else  
    .PMA_PLL0_REG_PLL_LOCKDET_REFCT           (6                             ),  
    .PMA_PLL0_REG_PLL_LOCKDET_FBCT            (6                             ),  
    .PMA_PLL0_REG_PLL_LOCKDET_ITER            (2                             ),
    `endif    
    .PMA_PLL0_REG_PLL_LOCKDET_LOCKCT          (4                             ),
    .PMA_PLL0_REG_PLL_UNLOCKDET_ITER          (2                             ),       
    .PMA_PLL0_REG_PD_VCO                      ("ON"                          ),                   
    .PMA_PLL0_REG_FBCLK_TEST_EN               ("FALSE"                       ),            
    .PMA_PLL0_REG_REFCLK_TEST_EN              ("FALSE"                       ),           
    .PMA_PLL0_REG_TEST_SEL                    (0                             ),                 
    .PMA_PLL0_REG_TEST_V_EN                   ("FALSE"                       ),                
    .PMA_PLL0_REG_TEST_SIG_HALF_EN            ("FALSE"                       ),         
    .PMA_PLL0_REG_TEST_FSM                    (0                             ),                   
    .PMA_PLL0_REG_REFCLK_OUT_PD               ("OFF"                         ), 
    .PMA_PLL0_REG_BGR_STARTUP_EN              ("FALSE"                       ),           
    .PMA_PLL0_REG_BGR_STARTUP                 ("FALSE"                       ),              
    .PMA_PLL0_REG_PD_BGR                      ("ON"                          ),                   
    .PMA_PLL0_REG_REFCLK_TERM_VCM_EN          ("TRUE"                        ),         
    .PMA_PLL0_REG_FBDIVA_5_EN                 ("TRUE"                        ), 
    .PMA_PLL0_REG_FBDIVB                      (2'b10                         ), 
    .PMA_PLL0_REG_RESET_N_PFDQP_OW            ("DISABLE"                     ),         
    .PMA_PLL0_REG_RESET_N_PFDQP               ("FALSE"                       ), 		           
    .PMA_PLL0_REG_QPCURRENT                   (4                             ),                
    .PMA_PLL0_REG_VC_FORCE_EN                 ("FALSE"                       ),              
    .PMA_PLL0_REG_VCRESET_C_RING              (4                             ),           
    .PMA_PLL0_REG_LPF_R_C                     (1                             ),                  
    .PMA_PLL0_REG_LPF_TR_C                    (0                             ),                 
    .PMA_PLL0_REG_PD_BIAS                     ("ON"                          ),                  
    .PMA_PLL0_REG_ICTRL_PLL                   (1                             ),                
    .PMA_PLL0_REG_BIAS_QP                     (1                             ),                  
    .PMA_PLL0_REG_BIAS_LANE_SYNC              (1                             ),           
    .PMA_PLL0_REG_BIAS_CLKBUFS1               (1                             ),             
    .PMA_PLL0_REG_TXPCLK_SEL                  (2                             ),               
    .PMA_PLL0_REG_BIAS_CLKBUFS3               (1                             ),            
    .PMA_PLL0_REG_LANE_SYNC_EN                ("TRUE"                        ),             
    .PMA_PLL0_REG_LANE_SYNC_EN_OW             ("ENABLE"                      ),          
    .PMA_PLL0_REG_BIAS_D2S                    (1                             ),                 
    .PMA_PLL0_REG_BIAS_REFD2S_C               (1                             ),            
    .PMA_PLL0_REG_BIAS_VCRST_C                (1                             ),             
    .PMA_PLL0_REG_BIAS_REFBUF_C               (1                             ),            
    .PMA_PLL0_REG_CLKBUFS1_C                  (1                             ),               
    .PMA_PLL0_REG_CLKBUFS2_C                  (6                             ),               
    .PMA_PLL0_REG_CLKBUFS3_C                  (6                             ),               
    .PMA_PLL0_REG_CLKBUFS4_C                  (1                             ),                 
    .PMA_PLL0_REG_PLL_REFCLK_CML_SEL          (0                             ), 
    .PMA_PLL0_REG_REFCLK_SEL                  ("FALSE"                       ), 
    .PMA_PLL0_REG_RESCAL_R_CODE_SIGN          ("TRUE"                        ),       
    .PMA_PLL0_REG_PLL_UNLOCKED_OW             ("DISABLE"                     ),          
    .PMA_PLL0_REG_PLL_UNLOCKED                ("FALSE"                       ),               
    .PMA_PLL0_REG_PLL_LOCKDET_MODE            ("FALSE"                       ), 
    .PMA_PLL0_REG_PLL_CLKBUF_PD_LEFT          ("ON"                          ), 
    .PMA_PLL0_REG_PLL_CLKBUF_PD_RIGHT         ("ON"                          ), 
    .PMA_PLL0_REG_RESCAL_EN                   ("FALSE"                       ),                
    .PMA_PLL0_REG_RESCAL_I_CODE_VAL           (0                             ),        
    .PMA_PLL0_REG_RESCAL_I_CODE_OW            (0                             ),         
    .PMA_PLL0_REG_RESCAL_ITER_VALID_SEL       (0                             ),    
    .PMA_PLL0_REG_RESCAL_WAIT_SEL             (0                             ),          
    .PMA_PLL0_REG_I_CTRL_MAX                  (45                            ),               
    .PMA_PLL0_REG_I_CTRL_MIN                  (19                            ),                 
    .PMA_PLL0_REG_RESERVED_167_160            (8'd0                          ), 
    .PMA_PLL0_REG_RESERVED_175_168            (0                             ),
    .PMA_PLL0_REG_RESERVED_183_176            (0                             ),
    .PMA_PLL0_REG_RESERVED_191_184            (0                             ),
    .PARM_CFG_HSST_RSTN                       ("TRUE"                        ),                      
    .PARM_PLL0_POWERUP                        ("ON"                          ), 
    .PARM_PLL0_RSTN                           ("TRUE"                        ),                          
    .PMA_PLL1_REG_PLL_POWERDOWN_OW            ("DISABLE"                     ), 
    .PMA_PLL1_REG_PLL_POWERDOWN               ("ON"                          ),            
    .PMA_PLL1_REG_PLL_RESET_N_OW              ("DISABLE"                     ),           
    .PMA_PLL1_REG_PLL_RESET_N                 ("TRUE"                        ),              
    .PMA_PLL1_REG_PLL_READY_OW                ("DISABLE"                     ),             
    .PMA_PLL1_REG_PLL_READY                   ("FALSE"                       ),                
    .PMA_PLL1_REG_LANE_SYNC_OW                ("DISABLE"                     ),             
    .PMA_PLL1_REG_LANE_SYNC                   ("FALSE"                       ),                
    .PMA_PLL1_REG_LOCKDET_REPEAT              ("DISABLE"                     ),           
    .PMA_PLL1_REG_RESCAL_I_CODE_PMA           ("DISABLE"                     ),        
    .PMA_PLL1_REG_RESCAL_RESET_N_OW           ("DISABLE"                     ),        
    .PMA_PLL1_REG_RESCAL_RESET_N              ("FALSE"                       ),           
    .PMA_PLL1_REG_RESCAL_DONE_OW              ("DISABLE"                     ),           
    .PMA_PLL1_REG_RESCAL_DONE                 ("FALSE"                       ),              
    .PMA_PLL1_REG_RESCAL_CODE_OW              ("DISABLE"                     ),           
    .PMA_PLL1_REG_LDO_VREF_SEL                (2                             ),             
    .PMA_PLL1_REG_BIAS_VCOREP_C               (1                             ),            
    .PMA_PLL1_REG_RESCAL_I_CODE               (32                            ),            
    .PMA_PLL1_REG_RESCAL_ONCHIP_SMALL_OW      ("DISABLE"                     ),  
    .PMA_PLL1_REG_RESCAL_ONCHIP_SMALL         (0                             ),      
    .PMA_PLL1_REG_JTAG_OE                     ("DISABLE"                     ),                  
    .PMA_PLL1_REG_JTAG_AC_MODE                ("DISABLE"                     ),             
    .PMA_PLL1_REG_JTAG_VHYSTSEL               (0                             ),            
    .PMA_PLL1_REG_PLL_LOCKDET_EN_OW           ("DISABLE"                     ),        
    .PMA_PLL1_REG_PLL_LOCKDET_EN              ("FALSE"                       ),           
    .PMA_PLL1_REG_PLL_LOCKDET_RESET_N_OW      ("DISABLE"                     ),   
    .PMA_PLL1_REG_PLL_LOCKDET_RESET_N         ("FALSE"                       ),      
    .PMA_PLL1_REG_PLL_LOCKED_OW               ("DISABLE"                     ),            
    .PMA_PLL1_REG_PLL_LOCKED                  ("FALSE"                       ),               
    .PMA_PLL1_REG_PLL_LOCKED_STICKY_CLEAR     ("FALSE"                       ),  
    .PMA_PLL1_REG_PLL_UNLOCKED_STICKY_CLEAR   ("FALSE"                       ),
    .PMA_PLL1_REG_NOFBCLK_STICKY_CLEAR        ("FALSE"                       ),
    `ifdef IPML_HSST_SPEEDUP_SIM
    .PMA_PLL1_REG_PLL_LOCKDET_REFCT           (4                             ),
    .PMA_PLL1_REG_PLL_LOCKDET_FBCT            (4                             ),
    .PMA_PLL1_REG_PLL_LOCKDET_ITER            (0                             ),
    `else 
    .PMA_PLL1_REG_PLL_LOCKDET_REFCT           (6                             ), 
    .PMA_PLL1_REG_PLL_LOCKDET_FBCT            (6                             ), 
    .PMA_PLL1_REG_PLL_LOCKDET_ITER            (2                             ),
    `endif    
    .PMA_PLL1_REG_PLL_LOCKDET_LOCKCT          (4                             ),
    .PMA_PLL1_REG_PLL_UNLOCKDET_ITER          (2                             ),       
    .PMA_PLL1_REG_PD_VCO                      ("ON"                          ),                   
    .PMA_PLL1_REG_FBCLK_TEST_EN               ("FALSE"                       ),            
    .PMA_PLL1_REG_REFCLK_TEST_EN              ("FALSE"                       ),           
    .PMA_PLL1_REG_TEST_SEL                    (0                             ),                 
    .PMA_PLL1_REG_TEST_V_EN                   ("FALSE"                       ),                
    .PMA_PLL1_REG_TEST_SIG_HALF_EN            ("FALSE"                       ),         
    .PMA_PLL1_REG_TEST_FSM                    (0                             ),                   
    .PMA_PLL1_REG_REFCLK_OUT_PD               ("OFF"                         ), 
    .PMA_PLL1_REG_BGR_STARTUP_EN              ("FALSE"                       ),           
    .PMA_PLL1_REG_BGR_STARTUP                 ("FALSE"                       ),              
    .PMA_PLL1_REG_PD_BGR                      ("ON"                          ),                   
    .PMA_PLL1_REG_REFCLK_TERM_VCM_EN          ("TRUE"                        ),         
    .PMA_PLL1_REG_FBDIVA_5_EN                 ("FALSE"                       ), 
    .PMA_PLL1_REG_FBDIVB                      (2'b01                         ), 
    .PMA_PLL1_REG_RESET_N_PFDQP_OW            ("DISABLE"                     ),         
    .PMA_PLL1_REG_RESET_N_PFDQP               ("FALSE"                       ),            
    .PMA_PLL1_REG_QPCURRENT                   (4                             ),                
    .PMA_PLL1_REG_VC_FORCE_EN                 ("FALSE"                       ),              
    .PMA_PLL1_REG_VCRESET_C_RING              (4                             ),           
    .PMA_PLL1_REG_LPF_R_C                     (1                             ),                  
    .PMA_PLL1_REG_LPF_TR_C                    (0                             ),                 
    .PMA_PLL1_REG_PD_BIAS                     ("ON"                          ),                  
    .PMA_PLL1_REG_ICTRL_PLL                   (1                             ),                
    .PMA_PLL1_REG_BIAS_QP                     (1                             ),                  
    .PMA_PLL1_REG_BIAS_LANE_SYNC              (1                             ),           
    .PMA_PLL1_REG_BIAS_CLKBUFS1               (1                             ),             
    .PMA_PLL1_REG_TXPCLK_SEL                  (0                             ),               
    .PMA_PLL1_REG_BIAS_CLKBUFS3               (1                             ),            
    .PMA_PLL1_REG_LANE_SYNC_EN                ("TRUE"                        ),             
    .PMA_PLL1_REG_LANE_SYNC_EN_OW             ("ENABLE"                      ),          
    .PMA_PLL1_REG_BIAS_D2S                    (1                             ),                 
    .PMA_PLL1_REG_BIAS_REFD2S_C               (1                             ),            
    .PMA_PLL1_REG_BIAS_VCRST_C                (1                             ),             
    .PMA_PLL1_REG_BIAS_REFBUF_C               (1                             ),            
    .PMA_PLL1_REG_CLKBUFS1_C                  (1                             ),               
    .PMA_PLL1_REG_CLKBUFS2_C                  (6                             ),               
    .PMA_PLL1_REG_CLKBUFS3_C                  (6                             ),               
    .PMA_PLL1_REG_CLKBUFS4_C                  (1                             ),                 
    .PMA_PLL1_REG_PLL_REFCLK_CML_SEL          (0                           ), 
    .PMA_PLL1_REG_REFCLK_SEL                  ("FALSE"                       ), 
    .PMA_PLL1_REG_RESCAL_R_CODE_SIGN          ("TRUE"                        ),       
    .PMA_PLL1_REG_PLL_UNLOCKED_OW             ("DISABLE"                     ),          
    .PMA_PLL1_REG_PLL_UNLOCKED                ("FALSE"                       ),               
    .PMA_PLL1_REG_PLL_LOCKDET_MODE            ("FALSE"                       ), 
    .PMA_PLL1_REG_PLL_CLKBUF_PD_LEFT          ("OFF"                         ), 
    .PMA_PLL1_REG_PLL_CLKBUF_PD_RIGHT         ("OFF"                         ), 
    .PMA_PLL1_REG_RESCAL_EN                   ("FALSE"                       ),                
    .PMA_PLL1_REG_RESCAL_I_CODE_VAL           (0                             ),        
    .PMA_PLL1_REG_RESCAL_I_CODE_OW            (0                             ),         
    .PMA_PLL1_REG_RESCAL_ITER_VALID_SEL       (0                             ),    
    .PMA_PLL1_REG_RESCAL_WAIT_SEL             (0                             ),          
    .PMA_PLL1_REG_I_CTRL_MAX                  (45                            ),               
    .PMA_PLL1_REG_I_CTRL_MIN                  (19                            ),                 
    .PMA_PLL1_REG_RESERVED_167_160            (8'd0                          ), 
    .PMA_PLL1_REG_RESERVED_175_168            (0                             ),
    .PMA_PLL1_REG_RESERVED_183_176            (0                             ),
    .PMA_PLL1_REG_RESERVED_191_184            (0                             ),  
    .PARM_PLL1_POWERUP                        ("OFF"                         ), 
    .PARM_PLL1_RSTN                           ("TRUE"                        ),                        
    .PARM_GRSN_DIS                            ("TRUE"                        ),                         
    .PARM_CFG_RSTN                            ("TRUE"                        )                         
) U_GTP_HSST(
    .P_REFCLKP_0                              (P_REFCLKP_0                                      ), 
    .P_REFCLKN_0                              (P_REFCLKN_0                                      ), 
    .P_PLL_TEST_0                             (P_PLL_TEST_0                                     ),
    .P_REFCLKP_1                              (P_REFCLKP_1                                      ),        
    .P_REFCLKN_1                              (P_REFCLKN_1                                      ),             
    .P_PLL_TEST_1                             (P_PLL_TEST_1                                     ),
    .P_RX_SDP0                                (P_RX_SDP0                                        ),        
    .P_RX_SDN0                                (P_RX_SDN0                                        ),           
    .P_TX_SDP0                                (P_TX_SDP0                                        ),   
    .P_TX_SDN0                                (P_TX_SDN0                                        ),   
    .P_RX_SDP1                                (P_RX_SDP1                                        ),                                   
    .P_RX_SDN1                                (P_RX_SDN1                                        ),           
    .P_TX_SDP1                                (P_TX_SDP1                                        ),   
    .P_TX_SDN1                                (P_TX_SDN1                                        ),           
    .P_RX_SDP2                                (P_RX_SDP2                                        ),                                   
    .P_RX_SDN2                                (P_RX_SDN2                                        ),           
    .P_TX_SDP2                                (P_TX_SDP2                                        ),   
    .P_TX_SDN2                                (P_TX_SDN2                                        ),     
    .P_RX_SDP3                                (P_RX_SDP3                                        ),                                   
    .P_RX_SDN3                                (P_RX_SDN3                                        ),           
    .P_TX_SDP3                                (P_TX_SDP3                                        ),   
    .P_TX_SDN3                                (P_TX_SDN3                                        ),     
    .P_RX0_CLK_FR_CORE                        (P_RX0_CLK_FR_CORE                                ),       
    .P_RX1_CLK_FR_CORE                        (P_RX1_CLK_FR_CORE                                ),         
    .P_RX2_CLK_FR_CORE                        (P_RX2_CLK_FR_CORE                                ),         
    .P_RX3_CLK_FR_CORE                        (P_RX3_CLK_FR_CORE                                ),         
    .P_RX0_CLK2_FR_CORE                       (P_RX0_CLK2_FR_CORE                               ), 
    .P_RX1_CLK2_FR_CORE                       (P_RX1_CLK2_FR_CORE                               ), 
    .P_RX2_CLK2_FR_CORE                       (P_RX2_CLK2_FR_CORE                               ), 
    .P_RX3_CLK2_FR_CORE                       (P_RX3_CLK2_FR_CORE                               ), 
    .P_TX0_CLK_FR_CORE                        (P_TX0_CLK_FR_CORE                                ),       
    .P_TX1_CLK_FR_CORE                        (P_TX1_CLK_FR_CORE                                ),         
    .P_TX2_CLK_FR_CORE                        (P_TX2_CLK_FR_CORE                                ),         
    .P_TX3_CLK_FR_CORE                        (P_TX3_CLK_FR_CORE                                ), 
    .P_TX0_CLK2_FR_CORE                       (P_TX0_CLK2_FR_CORE                               ), 
    .P_TX1_CLK2_FR_CORE                       (P_TX1_CLK2_FR_CORE                               ), 
    .P_TX2_CLK2_FR_CORE                       (P_TX2_CLK2_FR_CORE                               ), 
    .P_TX3_CLK2_FR_CORE                       (P_TX3_CLK2_FR_CORE                               ), 
    .P_HSST_RST                               (P_HSST_RST                                       ),
    .P_PCS_RX_RST_0                           (P_PCS_RX_RST_0                                   ),
    .P_PCS_RX_RST_1                           (P_PCS_RX_RST_1                                   ),        
    .P_PCS_RX_RST_2                           (P_PCS_RX_RST_2                                   ),
    .P_PCS_RX_RST_3                           (P_PCS_RX_RST_3                                   ),        
    .P_PCS_TX_RST_0                           (P_PCS_TX_RST_0                                   ),
    .P_PCS_TX_RST_1                           (P_PCS_TX_RST_1                                   ),        
    .P_PCS_TX_RST_2                           (P_PCS_TX_RST_2                                   ),        
    .P_PCS_TX_RST_3                           (P_PCS_TX_RST_3                                   ),
    .P_PCS_CB_RST_0                           (P_PCS_CB_RST_0                                   ), 
    .P_PCS_CB_RST_1                           (P_PCS_CB_RST_1                                   ), 
    .P_PCS_CB_RST_2                           (P_PCS_CB_RST_2                                   ), 
    .P_PCS_CB_RST_3                           (P_PCS_CB_RST_3                                   ), 
    .P_RXGEAR_SLIP_0                          (P_RXGEAR_SLIP_0                                  ), 
    .P_RXGEAR_SLIP_1                          (P_RXGEAR_SLIP_1                                  ), 
    .P_RXGEAR_SLIP_2                          (P_RXGEAR_SLIP_2                                  ), 
    .P_RXGEAR_SLIP_3                          (P_RXGEAR_SLIP_3                                  ), 
    .P_CFG_CLK                                (P_CFG_CLK                                        ),   
    .P_CFG_RST                                (P_CFG_RST                                        ),   
    .P_CFG_PSEL                               (P_CFG_PSEL                                       ), 
    .P_CFG_ENABLE                             (P_CFG_ENABLE                                     ),
    .P_CFG_WRITE                              (P_CFG_WRITE                                      ), 
    .P_CFG_ADDR                               (P_CFG_ADDR                                       ),  
    .P_CFG_WDATA                              (P_CFG_WDATA                                      ), 
    .P_TDATA_0                                (P_TDATA_0                                        ),
    .P_TDATA_1                                (P_TDATA_1                                        ),
    .P_TDATA_2                                (P_TDATA_2                                        ),
    .P_TDATA_3                                (P_TDATA_3                                        ),
    .P_PCS_WORD_ALIGN_EN                      (P_PCS_WORD_ALIGN_EN                              ), 
    .P_RX_POLARITY_INVERT                     (P_RX_POLARITY_INVERT                             ),
    .P_CEB_ADETECT_EN                         (P_CEB_ADETECT_EN                                 ),    
    .P_PCS_MCB_EXT_EN                         (P_PCS_MCB_EXT_EN                                 ),    
    .P_PCS_NEAREND_LOOP                       (P_PCS_NEAREND_LOOP                               ),  
    .P_PCS_FAREND_LOOP                        (P_PCS_FAREND_LOOP                                ),   
    .P_PMA_NEAREND_PLOOP                      (P_PMA_NEAREND_PLOOP                              ), 
    .P_PMA_NEAREND_SLOOP                      (P_PMA_NEAREND_SLOOP                              ), 
    .P_PMA_FAREND_PLOOP                       (P_PMA_FAREND_PLOOP                               ), 
    .P_CFG_READY                              (P_CFG_READY                                      ),         
    .P_CFG_RDATA                              (P_CFG_RDATA                                      ),         
    .P_CFG_INT                                (P_CFG_INT                                        ),           
    .P_PCS_RX_MCB_STATUS                      (P_PCS_RX_MCB_STATUS                              ), 
    .P_PCS_LSM_SYNCED                         (P_PCS_LSM_SYNCED                                 ),    
    .P_RDATA_0                                (P_RDATA_0                                        ),
    .P_RDATA_1                                (P_RDATA_1                                        ),
    .P_RDATA_2                                (P_RDATA_2                                        ),
    .P_RDATA_3                                (P_RDATA_3                                        ),
    .P_RCLK2FABRIC                            (P_RCLK2FABRIC                                    ),    
    .P_TCLK2FABRIC                            (P_TCLK2FABRIC                                    ),    
    .P_RESCAL_RST_I                           (P_RESCAL_RST_I                                   ),          
    .P_RESCAL_I_CODE_I                        (P_RESCAL_I_CODE_I                                ),   
    .P_RESCAL_I_CODE_O                        (P_RESCAL_I_CODE_O                                ),
    .P_REFCK2CORE_0                           (P_REFCK2CORE_0                                   ),         
    .P_PLL_REF_CLK_0                          (P_PLL_REF_CLK_0                                  ),        
    .P_PLL_RST_0                              (P_PLL_RST_0                                      ), 
    .P_PLLPOWERDOWN_0                         (P_PLLPOWERDOWN_0                                 ),
    .P_PLL_READY_0                            (P_PLL_READY_0                                    ),          
    .P_LANE_SYNC_0                            (P_LANE_SYNC_0                                    ),          
    .P_LANE_SYNC_EN_0                         (P_LANE_SYNC_EN_0                                 ),       
    .P_RATE_CHANGE_TCLK_ON_0                  (P_RATE_CHANGE_TCLK_ON_0                          ),
    .P_REFCK2CORE_1                           (P_REFCK2CORE_1                                   ),         
    .P_PLL_REF_CLK_1                          (P_PLL_REF_CLK_1                                  ),        
    .P_PLL_RST_1                              (P_PLL_RST_1                                      ),            
    .P_PLLPOWERDOWN_1                         (P_PLLPOWERDOWN_1                                 ),       
    .P_PLL_READY_1                            (P_PLL_READY_1                                    ),          
    .P_LANE_SYNC_1                            (P_LANE_SYNC_1                                    ),          
    .P_LANE_SYNC_EN_1                         (P_LANE_SYNC_EN_1                                 ),       
    .P_RATE_CHANGE_TCLK_ON_1                  (P_RATE_CHANGE_TCLK_ON_1                          ),
    .P_LANE_PD_0                              (P_LANE_PD_0                                      ),         
    .P_LANE_RST_0                             (P_LANE_RST_0                                     ),        
    .P_RX_LANE_PD_0                           (P_RX_LANE_PD_0                                   ),      
    .P_RX_PMA_RST_0                           (P_RX_PMA_RST_0                                   ),
    .P_CTLE_ADP_RST_0                         (P_CTLE_ADP_RST_0                                 ),     
    .P_RX_SIGDET_STATUS_0                     (P_RX_SIGDET_STATUS_0                             ),
    .P_RX_SATA_COMINIT_0                      (P_RX_SATA_COMINIT_0                              ), 
    .P_RX_SATA_COMWAKE_0                      (P_RX_SATA_COMWAKE_0                              ), 
    .P_RX_LS_DATA_0                           (P_RX_LS_DATA_0                                   ),      
    .P_RX_READY_0                             (P_RX_READY_0                                     ),        
    .P_TEST_STATUS_0                          (P_TEST_STATUS_0                                  ),     
    .P_TX_DEEMP_0                             (P_TX_DEEMP_0                                     ),        
    .P_TX_LS_DATA_0                           (P_TX_LS_DATA_0                                   ),      
    .P_TX_BEACON_EN_0                         (P_TX_BEACON_EN_0                                 ),    
    .P_TX_SWING_0                             (P_TX_SWING_0                                     ),        
    .P_TX_RXDET_REQ_0                         (P_TX_RXDET_REQ_0                                 ),    
    .P_TX_RATE_0                              (P_TX_RATE_0                                      ),         
    .P_TX_BUSWIDTH_0                          (P_TX_BUSWIDTH_0                                  ),     
    .P_TX_MARGIN_0                            (P_TX_MARGIN_0                                    ),       
    .P_TX_RXDET_STATUS_0                      (P_TX_RXDET_STATUS_0                              ), 
    .P_TX_PMA_RST_0                           (P_TX_PMA_RST_0                                   ),      
    .P_TX_LANE_PD_0                           (P_TX_LANE_PD_0                                   ),      
    .P_RX_RATE_0                              (P_RX_RATE_0                                      ),         
    .P_RX_BUSWIDTH_0                          (P_RX_BUSWIDTH_0                                  ),     
    .P_RX_HIGHZ_0                             (P_RX_HIGHZ_0                                     ),        
    .P_CA_ALIGN_RX                            (P_CA_ALIGN_RX                                    ),       
    .P_CA_ALIGN_TX                            (P_CA_ALIGN_TX                                    ),       
    .P_CIM_CLK_ALIGNER_RX0                    (P_CIM_CLK_ALIGNER_RX0                            ),
    .P_CIM_CLK_ALIGNER_TX0                    (P_CIM_CLK_ALIGNER_TX0                            ),
    .P_CIM_DYN_DLY_SEL_RX0                    (P_CIM_DYN_DLY_SEL_RX0                            ),
    .P_CIM_DYN_DLY_SEL_TX0                    (P_CIM_DYN_DLY_SEL_TX0                            ),
    .P_CIM_START_ALIGN_RX0                    (P_CIM_START_ALIGN_RX0                            ),
    .P_CIM_START_ALIGN_TX0                    (P_CIM_START_ALIGN_TX0                            ),
    .P_LANE_PD_1                              (P_LANE_PD_1                                      ),         
    .P_LANE_RST_1                             (P_LANE_RST_1                                     ),        
    .P_RX_LANE_PD_1                           (P_RX_LANE_PD_1                                   ),      
    .P_RX_PMA_RST_1                           (P_RX_PMA_RST_1                                   ),      
    .P_CTLE_ADP_RST_1                         (P_CTLE_ADP_RST_1                                 ),
    .P_RX_SIGDET_STATUS_1                     (P_RX_SIGDET_STATUS_1                             ),
    .P_RX_SATA_COMINIT_1                      (P_RX_SATA_COMINIT_1                              ), 
    .P_RX_SATA_COMWAKE_1                      (P_RX_SATA_COMWAKE_1                              ), 
    .P_RX_LS_DATA_1                           (P_RX_LS_DATA_1                                   ),      
    .P_RX_READY_1                             (P_RX_READY_1                                     ),        
    .P_TEST_STATUS_1                          (P_TEST_STATUS_1                                  ),     
    .P_TX_DEEMP_1                             (P_TX_DEEMP_1                                     ),        
    .P_TX_LS_DATA_1                           (P_TX_LS_DATA_1                                   ),      
    .P_TX_BEACON_EN_1                         (P_TX_BEACON_EN_1                                 ),    
    .P_TX_SWING_1                             (P_TX_SWING_1                                     ),        
    .P_TX_RXDET_REQ_1                         (P_TX_RXDET_REQ_1                                 ),    
    .P_TX_RATE_1                              (P_TX_RATE_1                                      ),         
    .P_TX_BUSWIDTH_1                          (P_TX_BUSWIDTH_1                                  ),     
    .P_TX_MARGIN_1                            (P_TX_MARGIN_1                                    ),       
    .P_TX_RXDET_STATUS_1                      (P_TX_RXDET_STATUS_1                              ), 
    .P_TX_PMA_RST_1                           (P_TX_PMA_RST_1                                   ),      
    .P_TX_LANE_PD_1                           (P_TX_LANE_PD_1                                   ),      
    .P_RX_RATE_1                              (P_RX_RATE_1                                      ),         
    .P_RX_BUSWIDTH_1                          (P_RX_BUSWIDTH_1                                  ),     
    .P_RX_HIGHZ_1                             (P_RX_HIGHZ_1                                     ),        
    .P_CIM_CLK_ALIGNER_RX1                    (P_CIM_CLK_ALIGNER_RX1                            ),
    .P_CIM_CLK_ALIGNER_TX1                    (P_CIM_CLK_ALIGNER_TX1                            ),
    .P_CIM_DYN_DLY_SEL_RX1                    (P_CIM_DYN_DLY_SEL_RX1                            ),
    .P_CIM_DYN_DLY_SEL_TX1                    (P_CIM_DYN_DLY_SEL_TX1                            ),
    .P_CIM_START_ALIGN_RX1                    (P_CIM_START_ALIGN_RX1                            ),
    .P_CIM_START_ALIGN_TX1                    (P_CIM_START_ALIGN_TX1                            ),
    .P_LANE_PD_2                              (P_LANE_PD_2                                      ),         
    .P_LANE_RST_2                             (P_LANE_RST_2                                     ),        
    .P_RX_LANE_PD_2                           (P_RX_LANE_PD_2                                   ),      
    .P_RX_PMA_RST_2                           (P_RX_PMA_RST_2                                   ),      
    .P_CTLE_ADP_RST_2                         (P_CTLE_ADP_RST_2                                 ),
    .P_RX_SIGDET_STATUS_2                     (P_RX_SIGDET_STATUS_2                             ),
    .P_RX_SATA_COMINIT_2                      (P_RX_SATA_COMINIT_2                              ), 
    .P_RX_SATA_COMWAKE_2                      (P_RX_SATA_COMWAKE_2                              ), 
    .P_RX_LS_DATA_2                           (P_RX_LS_DATA_2                                   ),      
    .P_RX_READY_2                             (P_RX_READY_2                                     ),        
    .P_TEST_STATUS_2                          (P_TEST_STATUS_2                                  ),     
    .P_TX_DEEMP_2                             (P_TX_DEEMP_2                                     ),        
    .P_TX_LS_DATA_2                           (P_TX_LS_DATA_2                                   ),      
    .P_TX_BEACON_EN_2                         (P_TX_BEACON_EN_2                                 ),    
    .P_TX_SWING_2                             (P_TX_SWING_2                                     ),        
    .P_TX_RXDET_REQ_2                         (P_TX_RXDET_REQ_2                                 ),    
    .P_TX_RATE_2                              (P_TX_RATE_2                                      ),         
    .P_TX_BUSWIDTH_2                          (P_TX_BUSWIDTH_2                                  ),     
    .P_TX_MARGIN_2                            (P_TX_MARGIN_2                                    ),       
    .P_TX_RXDET_STATUS_2                      (P_TX_RXDET_STATUS_2                              ), 
    .P_TX_PMA_RST_2                           (P_TX_PMA_RST_2                                   ),      
    .P_TX_LANE_PD_2                           (P_TX_LANE_PD_2                                   ),      
    .P_RX_RATE_2                              (P_RX_RATE_2                                      ),         
    .P_RX_BUSWIDTH_2                          (P_RX_BUSWIDTH_2                                  ),     
    .P_RX_HIGHZ_2                             (P_RX_HIGHZ_2                                     ),        
    .P_CIM_CLK_ALIGNER_RX2                    (P_CIM_CLK_ALIGNER_RX2                            ),
    .P_CIM_CLK_ALIGNER_TX2                    (P_CIM_CLK_ALIGNER_TX2                            ),
    .P_CIM_DYN_DLY_SEL_RX2                    (P_CIM_DYN_DLY_SEL_RX2                            ),
    .P_CIM_DYN_DLY_SEL_TX2                    (P_CIM_DYN_DLY_SEL_TX2                            ),
    .P_CIM_START_ALIGN_RX2                    (P_CIM_START_ALIGN_RX2                            ),
    .P_CIM_START_ALIGN_TX2                    (P_CIM_START_ALIGN_TX2                            ),
    .P_LANE_PD_3                              (P_LANE_PD_3                                      ),         
    .P_LANE_RST_3                             (P_LANE_RST_3                                     ),        
    .P_RX_LANE_PD_3                           (P_RX_LANE_PD_3                                   ),      
    .P_RX_PMA_RST_3                           (P_RX_PMA_RST_3                                   ),      
    .P_CTLE_ADP_RST_3                         (P_CTLE_ADP_RST_3                                 ),
    .P_RX_SIGDET_STATUS_3                     (P_RX_SIGDET_STATUS_3                             ),
    .P_RX_SATA_COMINIT_3                      (P_RX_SATA_COMINIT_3                              ), 
    .P_RX_SATA_COMWAKE_3                      (P_RX_SATA_COMWAKE_3                              ), 
    .P_RX_LS_DATA_3                           (P_RX_LS_DATA_3                                   ),      
    .P_RX_READY_3                             (P_RX_READY_3                                     ),        
    .P_TEST_STATUS_3                          (P_TEST_STATUS_3                                  ),     
    .P_TX_DEEMP_3                             (P_TX_DEEMP_3                                     ),        
    .P_TX_LS_DATA_3                           (P_TX_LS_DATA_3                                   ),      
    .P_TX_BEACON_EN_3                         (P_TX_BEACON_EN_3                                 ),    
    .P_TX_SWING_3                             (P_TX_SWING_3                                     ),        
    .P_TX_RXDET_REQ_3                         (P_TX_RXDET_REQ_3                                 ),    
    .P_TX_RATE_3                              (P_TX_RATE_3                                      ),         
    .P_TX_BUSWIDTH_3                          (P_TX_BUSWIDTH_3                                  ),     
    .P_TX_MARGIN_3                            (P_TX_MARGIN_3                                    ),       
    .P_TX_RXDET_STATUS_3                      (P_TX_RXDET_STATUS_3                              ), 
    .P_TX_PMA_RST_3                           (P_TX_PMA_RST_3                                   ),      
    .P_TX_LANE_PD_3                           (P_TX_LANE_PD_3                                   ),      
    .P_RX_RATE_3                              (P_RX_RATE_3                                      ),         
    .P_RX_BUSWIDTH_3                          (P_RX_BUSWIDTH_3                                  ),     
    .P_RX_HIGHZ_3                             (P_RX_HIGHZ_3                                     ),        
    .P_CIM_CLK_ALIGNER_RX3                    (P_CIM_CLK_ALIGNER_RX3                            ),
    .P_CIM_CLK_ALIGNER_TX3                    (P_CIM_CLK_ALIGNER_TX3                            ),
    .P_CIM_DYN_DLY_SEL_RX3                    (P_CIM_DYN_DLY_SEL_RX3                            ),
    .P_CIM_DYN_DLY_SEL_TX3                    (P_CIM_DYN_DLY_SEL_TX3                            ),
    .P_CIM_START_ALIGN_RX3                    (P_CIM_START_ALIGN_RX3                            ),
    .P_CIM_START_ALIGN_TX3                    (P_CIM_START_ALIGN_TX3                            ) 
);

endmodule
