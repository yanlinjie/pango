version https://git-lfs.github.com/spec/v1
oid sha256:fcb84b35e06b5557a2cef6d3f3a78e05aef34d12b0f63aa6d000ff4351df3658
size 5023
