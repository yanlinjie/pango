version https://git-lfs.github.com/spec/v1
oid sha256:37dcbd86e16bb3137437a9297e9af693cd01e04590e4413d02d142a7311a8db9
size 694
