version https://git-lfs.github.com/spec/v1
oid sha256:25043d69979aad94d19d7a146be9bea3fce15d8c3821e33b44087d3faad7d779
size 4458
